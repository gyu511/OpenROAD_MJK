VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "|" ;

PROPERTYDEFINITIONS
END PROPERTYDEFINITIONS

UNITS
    DATABASE MICRONS 2000 ;
END UNITS
SITE CoreSiteDie1
    CLASS CORE ;
    SIZE 0.141 BY 1.209 ;
END CoreSiteDie1

LAYER Metal1Die1
    TYPE ROUTING ;
    PITCH 0.19 ;
    WIDTH 0.06 ;
    AREA 0.02 ;
    SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025  ;
SPACINGTABLE
  PARALLELRUNLENGTH 0.000
  WIDTH 0.000	 0.060
  WIDTH 0.100	 0.100
  WIDTH 0.750	 0.250
  WIDTH 1.500	 0.450 ;
    DIRECTION HORIZONTAL ;
END Metal1Die1

MACRO OAI2BB1X4
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1135 0.82 1.156 1.018 ;
              RECT  0.042 0.82 1.156 0.8625 ;
              RECT  0.774 0.403 0.9615 0.445 ;
              RECT  0.8235 0.82 0.866 1.018 ;
              RECT  0.081 0.417 0.8095 0.4595 ;
              RECT  0.5265 0.82 0.569 1.018 ;
              RECT  0.3605 0.403 0.445 0.4595 ;
              RECT  0.2365 0.82 0.279 1.018 ;
              RECT  0.042 0.6925 0.1235 0.8625 ;
              RECT  0.081 0.417 0.1235 0.8625 ;
        END
    END Y
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3325 0.5795 1.4845 0.636 ;
              RECT  1.3325 0.4415 1.389 0.636 ;
              RECT  1.269 0.4415 1.389 0.4985 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.6925 1.796 0.82 ;
              RECT  1.6685 0.6925 1.796 0.7495 ;
              RECT  1.6685 0.537 1.725 0.7495 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.194 0.53 1.1985 0.5725 ;
              RECT  0.325 0.53 0.3815 0.6505 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END OAI2BB1X4

MACRO OA22X2
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.403 1.1415 0.445 ;
              RECT  1.032 0.403 1.0885 0.516 ;
              RECT  1.018 0.4735 1.0605 0.986 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.6925 0.9475 0.7845 ;
              RECT  0.707 0.6925 0.9475 0.7495 ;
              RECT  0.707 0.6925 0.7635 0.827 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.477 0.3815 0.8305 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.477 0.24 0.8305 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.477 0.523 0.8305 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END OA22X2

MACRO NAND3X8
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1995 0.6925 3.27 1.032 ;
              RECT  3.2275 0.286 3.27 1.032 ;
              RECT  0.548 0.286 3.27 0.3285 ;
              RECT  2.9095 0.742 3.27 0.7845 ;
              RECT  3.1535 0.6925 3.27 0.7845 ;
              RECT  2.9095 0.7175 2.952 1.032 ;
              RECT  0.2225 0.8555 2.952 0.898 ;
              RECT  2.6195 0.7495 2.662 1.032 ;
              RECT  2.305 0.8555 2.3475 0.94 ;
              RECT  2.015 0.8555 2.0575 0.94 ;
              RECT  1.725 0.8555 1.7675 0.94 ;
              RECT  1.4315 0.8555 1.474 0.94 ;
              RECT  1.117 0.7495 1.1595 1.032 ;
              RECT  0.827 0.8555 0.8695 0.94 ;
              RECT  0.537 0.8555 0.5795 0.94 ;
              RECT  0.2225 0.8445 0.265 1.032 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.6375 0.6255 2.729 0.668 ;
              RECT  2.5065 0.636 2.6795 0.6785 ;
              RECT  1.23 0.742 2.549 0.7845 ;
              RECT  2.5065 0.636 2.549 0.7845 ;
              RECT  1.8455 0.6255 1.8875 0.7845 ;
              RECT  1.803 0.6255 1.8875 0.668 ;
              RECT  1.23 0.636 1.2725 0.7845 ;
              RECT  0.905 0.636 1.2725 0.6785 ;
              RECT  0.905 0.6255 0.9895 0.6785 ;
              RECT  0.3355 0.742 0.9475 0.7845 ;
              RECT  0.905 0.6255 0.9475 0.7845 ;
              RECT  0.1975 0.7315 0.378 0.774 ;
              RECT  0.1975 0.5585 0.24 0.774 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.853 0.5125 3.0015 0.6325 ;
              RECT  2.4815 0.5125 3.0015 0.555 ;
              RECT  2.3935 0.523 2.5665 0.5655 ;
              RECT  2.1 0.629 2.4355 0.6715 ;
              RECT  2.3935 0.523 2.4355 0.6715 ;
              RECT  2.1 0.523 2.1425 0.6715 ;
              RECT  1.9585 0.523 2.1425 0.5655 ;
              RECT  1.6545 0.5125 2.001 0.555 ;
              RECT  1.612 0.523 1.697 0.5655 ;
              RECT  1.3435 0.629 1.6545 0.6715 ;
              RECT  1.612 0.523 1.6545 0.6715 ;
              RECT  1.3435 0.523 1.3855 0.6715 ;
              RECT  1.0605 0.523 1.3855 0.5655 ;
              RECT  0.735 0.5125 1.103 0.555 ;
              RECT  0.449 0.629 0.7775 0.6715 ;
              RECT  0.735 0.5125 0.7775 0.6715 ;
              RECT  0.318 0.6185 0.491 0.661 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.072 0.523 3.157 0.5655 ;
              RECT  3.072 0.3995 3.1145 0.5655 ;
              RECT  0.622 0.3995 3.1145 0.4415 ;
              RECT  2.2375 0.516 2.3225 0.5585 ;
              RECT  2.28 0.3995 2.3225 0.5585 ;
              RECT  1.4565 0.516 1.541 0.5585 ;
              RECT  1.4565 0.3995 1.499 0.5585 ;
              RECT  0.562 0.516 0.6645 0.5585 ;
              RECT  0.608 0.424 0.6645 0.5585 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END NAND3X8

MACRO SDFFRX4
    CLASS CORE ;
    SIZE 5.515 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.6665 0.3425 5.084 0.385 ;
              RECT  5.0275 0.6715 5.0695 0.9475 ;
              RECT  4.709 0.6715 5.0695 0.714 ;
              RECT  4.709 0.6715 4.78 0.9475 ;
              RECT  4.709 0.5585 4.7655 0.9475 ;
              RECT  4.709 0.3425 4.7515 0.9475 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4475 0.6715 4.49 0.9475 ;
              RECT  4.1435 0.6715 4.49 0.714 ;
              RECT  4.002 0.3425 4.419 0.385 ;
              RECT  4.1435 0.5585 4.2 0.9475 ;
              RECT  4.1435 0.3425 4.186 0.9475 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.783 0.4525 3.825 0.537 ;
              RECT  3.2985 0.456 3.825 0.4985 ;
              RECT  3.341 0.4525 3.825 0.4985 ;
              RECT  3.341 0.2755 3.3835 0.4985 ;
              RECT  3.118 0.2755 3.3835 0.318 ;
              RECT  3.118 0.2085 3.1605 0.318 ;
              RECT  2.6195 0.2085 3.1605 0.251 ;
              RECT  2.28 0.569 2.662 0.6115 ;
              RECT  2.6195 0.2085 2.662 0.6115 ;
              RECT  2.57 0.4415 2.662 0.4985 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.424 1.0885 0.7775 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.424 0.9475 0.7775 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.4805 0.7775 ;
              RECT  0.325 0.523 0.3815 0.7775 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7775 0.18 0.82 0.7775 ;
              RECT  0.3815 0.18 0.82 0.2225 ;
              RECT  0.449 0.4415 0.5335 0.484 ;
              RECT  0.1975 0.41 0.491 0.4525 ;
              RECT  0.3815 0.18 0.424 0.4525 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.515 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.515 0.042 ;
        END
    END VSS
END SDFFRX4

MACRO TLATSRX1
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.622 0.2895 0.6645 0.7565 ;
              RECT  0.608 0.424 0.6645 0.516 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.159 0.2895 0.2155 0.912 ;
              RECT  0.042 0.2895 0.2155 0.3815 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.5975 2.4535 0.8165 ;
              RECT  2.397 0.555 2.4535 0.8165 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4315 0.576 1.718 0.6785 ;
              RECT  1.4315 0.555 1.488 0.6785 ;
        END
    END RN
    PIN G
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.131 0.576 1.248 0.6325 ;
              RECT  1.131 0.576 1.1875 0.8695 ;
        END
    END G
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.4595 0.9475 0.7705 ;
              RECT  0.8485 0.5935 0.9475 0.6505 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END TLATSRX1

MACRO OAI2BB1X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.5585 0.24 0.9475 ;
              RECT  0.0845 0.5585 0.24 0.601 ;
              RECT  0.0845 0.2825 0.127 0.601 ;
              RECT  0.042 0.2895 0.127 0.3815 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.3815 0.7915 ;
              RECT  0.311 0.4525 0.3675 0.7495 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4525 0.5515 0.523 0.7915 ;
              RECT  0.4525 0.4525 0.509 0.7915 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6925 0.806 0.7845 ;
              RECT  0.707 0.4735 0.7635 0.7495 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OAI2BB1X1

MACRO DLY4X1
    CLASS CORE ;
    SIZE 4.101 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.4415 0.3995 0.4985 ;
              RECT  0.3075 0.3815 0.364 0.912 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.8605 0.4875 3.917 0.841 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.101 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.101 0.042 ;
        END
    END VSS
END DLY4X1

MACRO ADDFX4
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.6945 0.424 3.7755 0.516 ;
              RECT  3.355 0.707 3.737 0.7495 ;
              RECT  3.6945 0.35 3.737 0.7495 ;
              RECT  3.652 0.293 3.6945 0.392 ;
              RECT  3.645 0.707 3.6875 0.9825 ;
              RECT  3.355 0.35 3.737 0.392 ;
              RECT  3.355 0.707 3.3975 0.9825 ;
              RECT  3.355 0.293 3.3975 0.392 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.537 0.6505 0.5795 0.9155 ;
              RECT  0.1835 0.424 0.5795 0.4665 ;
              RECT  0.537 0.3675 0.5795 0.4665 ;
              RECT  0.1975 0.6505 0.5795 0.6925 ;
              RECT  0.24 0.6505 0.2825 0.9155 ;
              RECT  0.24 0.3675 0.2825 0.4665 ;
              RECT  0.1975 0.424 0.24 0.6925 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.245 0.5795 3.058 0.622 ;
              RECT  1.598 0.622 2.287 0.6645 ;
              RECT  1.598 0.5585 1.785 0.6645 ;
              RECT  1.248 0.5585 1.785 0.601 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1285 0.4415 3.171 0.5265 ;
              RECT  2.9945 0.4415 3.171 0.509 ;
              RECT  2.1315 0.4665 3.171 0.509 ;
              RECT  1.856 0.509 2.174 0.5515 ;
              RECT  1.856 0.445 1.8985 0.5515 ;
              RECT  1.0885 0.445 1.8985 0.4875 ;
              RECT  1.0885 0.445 1.131 0.53 ;
        END
    END A
    PIN CI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.955 0.3535 2.839 0.3955 ;
              RECT  1.976 0.3535 2.061 0.438 ;
              RECT  1.58 0.332 1.9975 0.3745 ;
              RECT  1.58 0.3075 1.672 0.3745 ;
        END
    END CI
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END ADDFX4

MACRO CLKAND2X12
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.853 0.647 2.927 0.9685 ;
              RECT  2.8705 0.5585 2.927 0.9685 ;
              RECT  2.8705 0.4205 2.913 0.9685 ;
              RECT  1.6295 0.4205 2.913 0.463 ;
              RECT  1.6935 0.647 2.927 0.689 ;
              RECT  2.7895 0.247 2.8315 0.463 ;
              RECT  2.563 0.647 2.6055 0.9685 ;
              RECT  2.4995 0.247 2.542 0.463 ;
              RECT  2.273 0.647 2.3155 0.9685 ;
              RECT  2.2095 0.247 2.252 0.463 ;
              RECT  1.983 0.647 2.0255 0.9685 ;
              RECT  1.9195 0.247 1.962 0.463 ;
              RECT  1.6935 0.647 1.7355 0.9685 ;
              RECT  1.6295 0.247 1.672 0.463 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2975 0.576 1.446 0.6185 ;
              RECT  0.4665 0.6715 1.389 0.714 ;
              RECT  1.2975 0.576 1.389 0.714 ;
              RECT  0.841 0.629 0.8835 0.714 ;
              RECT  0.4665 0.629 0.509 0.714 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.117 0.516 1.1595 0.601 ;
              RECT  0.339 0.516 1.1595 0.5585 ;
              RECT  0.682 0.516 0.767 0.5655 ;
              RECT  0.325 0.5585 0.3815 0.6505 ;
              RECT  0.187 0.5585 0.3815 0.601 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END CLKAND2X12

MACRO MXI3XL
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.3675 2.3615 0.721 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.061 0.5585 2.227 0.767 ;
              RECT  2.061 0.523 2.1175 0.767 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.6645 1.8135 0.721 ;
              RECT  1.4385 0.576 1.5305 0.721 ;
        END
    END S1
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.951 0.5975 1.0885 0.8025 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3005 0.576 0.654 0.6325 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.7035 0.636 0.76 ;
              RECT  0.166 0.7105 0.258 0.767 ;
              RECT  0.173 0.682 0.2295 0.767 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END MXI3XL

MACRO NAND3X6
    CLASS CORE ;
    SIZE 2.9695 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2755 0.834 2.927 0.8765 ;
              RECT  2.8845 0.3815 2.927 0.8765 ;
              RECT  2.8705 0.6925 2.927 0.8765 ;
              RECT  2.4075 0.3815 2.927 0.424 ;
              RECT  2.7115 0.834 2.754 1.011 ;
              RECT  2.4215 0.834 2.464 0.919 ;
              RECT  2.4075 0.226 2.45 0.424 ;
              RECT  1.389 0.304 2.45 0.346 ;
              RECT  2.1315 0.834 2.174 0.919 ;
              RECT  1.842 0.7565 1.884 1.011 ;
              RECT  1.534 0.834 1.5765 0.919 ;
              RECT  1.389 0.226 1.4315 0.424 ;
              RECT  0.548 0.226 1.4315 0.2685 ;
              RECT  1.1455 0.834 1.1875 0.919 ;
              RECT  0.8555 0.834 0.898 0.919 ;
              RECT  0.5655 0.834 0.608 0.919 ;
              RECT  0.548 0.226 0.59 0.424 ;
              RECT  0.2755 0.834 0.318 0.919 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7575 0.537 2.807 0.622 ;
              RECT  2.068 0.721 2.8 0.7635 ;
              RECT  2.7575 0.537 2.8 0.7635 ;
              RECT  2.068 0.643 2.1105 0.7635 ;
              RECT  1.7285 0.643 2.1105 0.6855 ;
              RECT  0.2435 0.721 1.771 0.7635 ;
              RECT  1.7285 0.643 1.771 0.7635 ;
              RECT  1.0075 0.643 1.092 0.7635 ;
              RECT  0.2435 0.576 0.286 0.7635 ;
              RECT  0.166 0.576 0.286 0.6325 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.181 0.608 2.683 0.6505 ;
              RECT  2.588 0.5585 2.6445 0.6505 ;
              RECT  2.181 0.53 2.2235 0.6505 ;
              RECT  1.6155 0.53 2.2235 0.5725 ;
              RECT  1.163 0.608 1.658 0.6505 ;
              RECT  1.6155 0.53 1.658 0.6505 ;
              RECT  1.163 0.53 1.2055 0.6505 ;
              RECT  0.894 0.53 1.2055 0.5725 ;
              RECT  0.781 0.569 0.9365 0.6115 ;
              RECT  0.357 0.608 0.8235 0.6505 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.2945 0.4945 2.4145 0.537 ;
              RECT  2.2945 0.417 2.3365 0.537 ;
              RECT  1.5025 0.417 2.3365 0.4595 ;
              RECT  1.276 0.4945 1.545 0.537 ;
              RECT  1.5025 0.417 1.545 0.537 ;
              RECT  1.276 0.417 1.3185 0.537 ;
              RECT  0.781 0.417 1.3185 0.4595 ;
              RECT  0.668 0.4415 0.8235 0.4985 ;
              RECT  0.6255 0.4945 0.7105 0.537 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.9695 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.9695 0.042 ;
        END
    END VSS
END NAND3X6

MACRO SDFFRX2
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7455 0.643 0.8305 0.7 ;
              RECT  0.7455 0.424 0.806 0.516 ;
              RECT  0.7455 0.346 0.8025 0.7 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4595 0.424 0.523 0.516 ;
              RECT  0.3955 0.643 0.516 0.7 ;
              RECT  0.4595 0.346 0.516 0.7 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.285 0.424 4.3415 0.516 ;
              RECT  3.9845 0.424 4.3415 0.4805 ;
              RECT  3.9845 0.424 4.041 0.622 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1115 0.5515 4.1965 0.608 ;
              RECT  3.9845 0.7105 4.168 0.767 ;
              RECT  4.1115 0.5515 4.168 0.767 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.6305 0.424 3.6875 0.615 ;
              RECT  3.5775 0.5585 3.6345 0.7245 ;
        END
    END SI
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.9655 0.9755 2.6655 1.018 ;
              RECT  1.9655 0.742 2.008 1.018 ;
              RECT  1.739 0.742 2.008 0.7845 ;
              RECT  1.739 0.6925 1.796 0.7845 ;
              RECT  1.739 0.5935 1.7815 0.7845 ;
              RECT  1.686 0.5935 1.7815 0.636 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0145 0.403 1.1595 0.4985 ;
              RECT  1.0145 0.403 1.071 0.668 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END SDFFRX2

MACRO MX3X1
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0915 0.5405 0.134 0.951 ;
              RECT  0.0915 0.272 0.134 0.357 ;
              RECT  0.0565 0.2895 0.0985 0.583 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4705 0.7105 1.955 0.767 ;
              RECT  1.4705 0.682 1.527 0.767 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.548 1.916 0.6045 ;
              RECT  1.598 0.548 1.6545 0.6395 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.117 0.4595 1.1735 0.6925 ;
              RECT  1.032 0.4595 1.1735 0.516 ;
              RECT  1.032 0.424 1.0885 0.516 ;
        END
    END B
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.339 0.9475 0.6925 ;
        END
    END S1
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.4415 0.3815 0.795 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END MX3X1

MACRO SDFFSRHQX1
    CLASS CORE ;
    SIZE 5.515 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0775 0.4735 0.12 0.912 ;
              RECT  0.042 0.424 0.0985 0.516 ;
              RECT  0.0565 0.3605 0.0985 0.516 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.826 0.456 5.349 0.4985 ;
              RECT  5.2255 0.4415 5.349 0.4985 ;
              RECT  4.826 0.456 4.868 0.6395 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.0945 0.576 5.381 0.6325 ;
              RECT  5.0945 0.5725 5.19 0.6925 ;
              RECT  5.1155 0.569 5.19 0.6925 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.55 0.3815 4.642 0.643 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1365 0.576 4.4795 0.6325 ;
              RECT  4.1365 0.576 4.359 0.643 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.531 0.9365 3.026 0.979 ;
              RECT  2.531 0.82 2.5735 0.979 ;
              RECT  2.2625 0.82 2.5735 0.8625 ;
              RECT  1.697 0.9155 2.305 0.958 ;
              RECT  2.2625 0.82 2.305 0.958 ;
              RECT  1.697 0.668 1.739 0.958 ;
              RECT  1.0465 0.668 1.739 0.7105 ;
              RECT  1.0465 0.5585 1.0885 0.7105 ;
              RECT  1.032 0.5585 1.0885 0.6505 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.5585 0.9475 0.6505 ;
              RECT  0.7245 0.5585 0.9475 0.643 ;
              RECT  0.7245 0.463 0.781 0.643 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.515 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.515 0.042 ;
        END
    END VSS
END SDFFSRHQX1

MACRO TLATNTSCAX16
    CLASS CORE ;
    SIZE 5.374 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.0345 0.576 5.077 0.993 ;
              RECT  5.0025 0.371 5.045 0.6185 ;
              RECT  3.295 0.576 5.077 0.6185 ;
              RECT  4.7445 0.4135 5.045 0.456 ;
              RECT  4.7445 0.576 4.787 0.993 ;
              RECT  4.6915 0.403 4.7765 0.445 ;
              RECT  4.4545 0.576 4.497 0.993 ;
              RECT  4.4225 0.371 4.465 0.6185 ;
              RECT  4.1645 0.4135 4.465 0.456 ;
              RECT  4.1645 0.576 4.207 0.993 ;
              RECT  4.1115 0.403 4.1965 0.445 ;
              RECT  3.8745 0.576 3.917 0.993 ;
              RECT  3.843 0.371 3.8855 0.6185 ;
              RECT  3.585 0.4135 3.8855 0.456 ;
              RECT  3.585 0.576 3.627 0.993 ;
              RECT  3.5315 0.403 3.6165 0.445 ;
              RECT  3.295 0.5585 3.3515 0.6505 ;
              RECT  3.295 0.3955 3.3375 0.993 ;
              RECT  3.263 0.3535 3.3055 0.438 ;
        END
    END ECK
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.318 0.523 0.6715 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.318 0.3815 0.6715 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.3815 0.0985 0.6715 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.374 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.374 0.042 ;
        END
    END VSS
END TLATNTSCAX16

MACRO OAI33XL
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.682 0.8375 1.23 0.88 ;
              RECT  1.1875 0.1835 1.23 0.88 ;
              RECT  1.1735 0.6925 1.23 0.88 ;
              RECT  0.8485 0.3005 1.23 0.3425 ;
              RECT  1.1275 0.1835 1.23 0.3425 ;
              RECT  0.8485 0.205 0.8905 0.3425 ;
              RECT  0.806 0.205 0.8905 0.247 ;
              RECT  0.682 0.8375 0.7245 0.9685 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5265 0.3815 0.88 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.7105 0.799 0.767 ;
              RECT  0.608 0.548 0.6645 0.767 ;
        END
    END B2
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1555 0.4595 0.226 0.6505 ;
              RECT  0.042 0.4595 0.226 0.516 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END A0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5585 0.523 0.912 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.4135 0.9475 0.767 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.424 1.0885 0.753 ;
              RECT  1.018 0.4135 1.0745 0.4985 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OAI33XL

MACRO TLATSRX4
    CLASS CORE ;
    SIZE 5.374 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.899 0.477 3.125 0.5195 ;
              RECT  3.0825 0.3285 3.125 0.5195 ;
              RECT  2.5455 0.7035 2.9835 0.7455 ;
              RECT  2.899 0.477 2.9415 0.7455 ;
              RECT  2.588 0.5585 2.6445 0.7455 ;
              RECT  2.588 0.3285 2.63 0.7455 ;
        END
    END QN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.376 0.576 3.903 0.6325 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.041 0.219 4.1255 0.2615 ;
              RECT  3.772 0.247 4.0835 0.2895 ;
              RECT  3.4645 0.2155 3.8145 0.258 ;
              RECT  3.196 0.35 3.507 0.392 ;
              RECT  3.4645 0.2155 3.507 0.392 ;
              RECT  3.196 0.2155 3.2385 0.392 ;
              RECT  2.9695 0.2155 3.2385 0.258 ;
              RECT  2.701 0.364 3.012 0.4065 ;
              RECT  2.9695 0.2155 3.012 0.4065 ;
              RECT  2.701 0.2155 2.7435 0.4065 ;
              RECT  2.4745 0.2155 2.7435 0.258 ;
              RECT  2.2485 0.385 2.517 0.4275 ;
              RECT  2.4745 0.2155 2.517 0.4275 ;
              RECT  2.2485 0.2155 2.291 0.4275 ;
              RECT  2.022 0.2155 2.291 0.258 ;
              RECT  1.796 0.385 2.0645 0.4275 ;
              RECT  2.022 0.2155 2.0645 0.4275 ;
              RECT  1.796 0.2155 1.838 0.4275 ;
              RECT  1.5695 0.2155 1.838 0.258 ;
              RECT  1.3435 0.385 1.612 0.4275 ;
              RECT  1.5695 0.2155 1.612 0.4275 ;
              RECT  1.3435 0.2155 1.3855 0.4275 ;
              RECT  1.117 0.2155 1.3855 0.258 ;
              RECT  0.8905 0.385 1.1595 0.4275 ;
              RECT  1.117 0.2155 1.1595 0.4275 ;
              RECT  0.8905 0.2155 0.933 0.4275 ;
              RECT  0.6645 0.2155 0.933 0.258 ;
              RECT  0.4665 0.424 0.707 0.4665 ;
              RECT  0.6645 0.2155 0.707 0.4665 ;
              RECT  0.4665 0.424 0.523 0.516 ;
              RECT  0.4665 0.424 0.5195 0.5515 ;
        END
    END RN
    PIN G
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.021 0.562 0.2825 0.6325 ;
              RECT  0.1975 0.484 0.2825 0.6325 ;
        END
    END G
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.992 0.5585 5.0485 0.6505 ;
              RECT  4.822 0.5585 5.0485 0.643 ;
              RECT  4.822 0.4665 4.879 0.643 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7565 0.7035 1.2725 0.7455 ;
              RECT  1.23 0.3285 1.2725 0.7455 ;
              RECT  0.7775 0.5585 0.9475 0.7455 ;
              RECT  0.7775 0.3285 0.82 0.7455 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.374 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.374 0.042 ;
        END
    END VSS
END TLATSRX4

MACRO DFFHQX4
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.899 0.576 3.2525 0.6325 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.304 0.24 0.6575 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7705 0.6575 0.813 0.912 ;
              RECT  0.7385 0.3815 0.781 0.7 ;
              RECT  0.4665 0.4735 0.781 0.516 ;
              RECT  0.4805 0.403 0.523 0.912 ;
              RECT  0.4665 0.403 0.523 0.516 ;
              RECT  0.385 0.403 0.523 0.445 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END DFFHQX4

MACRO AOI221X2
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5695 0.7035 1.612 0.8025 ;
              RECT  0.7635 0.7035 1.612 0.7455 ;
              RECT  0.4275 0.318 1.534 0.3605 ;
              RECT  0.7635 0.318 0.806 0.7455 ;
              RECT  0.7495 0.5585 0.806 0.6505 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0145 0.576 1.368 0.6325 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5405 0.523 0.753 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2015 0.431 0.6785 0.4875 ;
              RECT  0.166 0.4415 0.258 0.5055 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.449 1.368 0.5055 ;
              RECT  1.156 0.4415 1.248 0.5055 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.46 0.576 1.8135 0.6325 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END AOI221X2

MACRO ADDFX2
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9875 0.728 3.072 0.7705 ;
              RECT  3.0085 0.424 3.0685 0.516 ;
              RECT  3.0085 0.2965 3.051 0.7705 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.194 0.3815 0.2365 0.926 ;
              RECT  0.042 0.5585 0.2365 0.601 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0075 0.5795 2.641 0.622 ;
              RECT  1.4565 0.5795 1.513 0.7845 ;
              RECT  0.841 0.5725 1.039 0.615 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7115 0.4665 2.8035 0.6325 ;
              RECT  1.0815 0.4665 2.8035 0.509 ;
              RECT  0.728 0.4595 1.11 0.502 ;
              RECT  0.6855 0.484 0.7705 0.5265 ;
        END
    END A
    PIN CI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.3535 2.485 0.3955 ;
              RECT  1.156 0.3075 1.248 0.3955 ;
        END
    END CI
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END ADDFX2

MACRO AOI22XL
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6395 0.788 0.682 0.873 ;
              RECT  0.636 0.608 0.6785 0.8305 ;
              RECT  0.4665 0.608 0.6785 0.6505 ;
              RECT  0.4665 0.5585 0.523 0.6505 ;
              RECT  0.4805 0.18 0.523 0.6505 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.318 0.24 0.6715 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.318 0.806 0.6715 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5935 0.424 0.6645 0.516 ;
              RECT  0.5935 0.1765 0.6505 0.516 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.205 0.3955 0.4945 ;
              RECT  0.325 0.1555 0.3815 0.247 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END AOI22XL

MACRO NAND3BX2
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8485 0.721 0.8905 0.951 ;
              RECT  0.2615 0.753 0.8905 0.795 ;
              RECT  0.5585 0.753 0.601 0.951 ;
              RECT  0.106 0.2365 0.583 0.279 ;
              RECT  0.2615 0.7105 0.304 0.951 ;
              RECT  0.106 0.7105 0.304 0.767 ;
              RECT  0.106 0.2365 0.148 0.767 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.622 0.576 0.6785 0.682 ;
              RECT  0.3745 0.576 0.6785 0.6325 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.5055 0.806 0.6505 ;
              RECT  0.332 0.463 0.799 0.5055 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0535 0.463 1.11 0.6505 ;
              RECT  1.032 0.555 1.0885 0.795 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END NAND3BX2

MACRO SDFFTRXL
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.318 0.721 0.403 ;
              RECT  0.608 0.318 0.6645 0.8555 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.159 0.3815 0.2155 0.721 ;
              RECT  0.042 0.424 0.2155 0.516 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.147 0.5125 4.391 0.569 ;
              RECT  4.267 0.403 4.391 0.569 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.864 0.4415 4.076 0.4985 ;
              RECT  3.864 0.4415 3.9205 0.6395 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.7015 0.4415 3.7935 0.76 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.906 0.364 2.9625 0.643 ;
              RECT  2.8705 0.5585 2.927 0.682 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8835 0.59 0.9685 0.647 ;
              RECT  0.735 0.7105 0.965 0.767 ;
              RECT  0.8835 0.59 0.965 0.767 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END SDFFTRXL

MACRO OR3X2
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7245 0.4735 0.9475 0.516 ;
              RECT  0.8905 0.424 0.9475 0.516 ;
              RECT  0.6575 0.643 0.767 0.6855 ;
              RECT  0.7245 0.2615 0.767 0.6855 ;
              RECT  0.6575 0.643 0.7 0.919 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4415 0.4415 0.5405 0.4985 ;
              RECT  0.4415 0.4415 0.5265 0.753 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2015 0.5585 0.258 0.7845 ;
              RECT  0.1835 0.449 0.24 0.6505 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.431 0.0985 0.7845 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END OR3X2

MACRO CLKBUFX2
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.247 0.6115 0.2895 0.933 ;
              RECT  0.247 0.35 0.2895 0.4345 ;
              RECT  0.2155 0.392 0.258 0.654 ;
              RECT  0.1835 0.424 0.258 0.516 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3605 0.7105 0.5405 0.767 ;
              RECT  0.484 0.537 0.5405 0.767 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END CLKBUFX2

MACRO TLATX1
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1705 0.3815 2.2375 0.9365 ;
              RECT  2.146 0.4415 2.2375 0.4985 ;
              RECT  2.153 0.3815 2.2375 0.4985 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.612 0.3815 1.6545 1.0005 ;
              RECT  1.598 0.424 1.6545 0.516 ;
        END
    END QN
    PIN G
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.5515 1.3715 0.905 ;
        END
    END G
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5125 0.449 0.7245 ;
              RECT  0.325 0.438 0.3815 0.7245 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END TLATX1

MACRO DFFHQX2
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.344 0.3815 2.386 0.6925 ;
              RECT  2.319 0.6505 2.3615 1.0355 ;
              RECT  2.305 0.6925 2.3615 0.7845 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5265 0.569 0.7385 0.6255 ;
              RECT  0.5265 0.569 0.682 0.767 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1445 0.4595 0.2015 0.6325 ;
              RECT  0.042 0.4595 0.2015 0.516 ;
              RECT  0.042 0.3815 0.0985 0.516 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END DFFHQX2

MACRO MXI4XL
    CLASS CORE ;
    SIZE 2.9695 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.095 0.3815 0.152 0.721 ;
              RECT  0.042 0.424 0.152 0.516 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4285 0.576 2.782 0.6325 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.464 0.7035 2.7505 0.7915 ;
              RECT  2.4285 0.7035 2.7505 0.767 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.962 0.7105 2.1315 0.767 ;
              RECT  1.962 0.5265 2.0185 0.767 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.626 0.622 1.8915 0.6785 ;
              RECT  1.626 0.622 1.8135 0.767 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.191 0.6395 1.2865 0.6965 ;
              RECT  1.191 0.4415 1.248 0.6965 ;
              RECT  1.131 0.4415 1.248 0.4985 ;
        END
    END D
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.94 0.1905 0.9825 0.6785 ;
              RECT  0.339 0.1905 0.9825 0.233 ;
              RECT  0.7495 0.173 0.834 0.233 ;
              RECT  0.339 0.502 0.385 0.5865 ;
              RECT  0.339 0.1905 0.3815 0.5865 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END S1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.9695 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.9695 0.042 ;
        END
    END VSS
END MXI4XL

MACRO AOI2BB2X2
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7745 0.7035 1.817 0.8025 ;
              RECT  1.329 0.7035 1.817 0.7455 ;
              RECT  1.6085 0.3145 1.6935 0.357 ;
              RECT  1.138 0.3285 1.651 0.371 ;
              RECT  1.4845 0.7035 1.527 0.8025 ;
              RECT  1.329 0.3285 1.3715 0.7455 ;
              RECT  1.315 0.5585 1.3715 0.6505 ;
              RECT  0.993 0.3145 1.1805 0.357 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.467 0.569 1.8135 0.6325 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.442 0.4415 1.8595 0.4985 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.424 0.3815 0.7775 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.325 0.24 0.6785 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END AOI2BB2X2

MACRO SEDFFTRX2
    CLASS CORE ;
    SIZE 5.798 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5245 0.3675 3.6695 0.424 ;
              RECT  3.5245 0.3675 3.581 0.721 ;
              RECT  3.4365 0.424 3.581 0.516 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.2525 0.5585 3.3515 0.6505 ;
              RECT  3.2525 0.3675 3.3375 0.424 ;
              RECT  3.2065 0.6255 3.3125 0.7 ;
              RECT  3.2525 0.3675 3.309 0.7 ;
              RECT  3.2065 0.6255 3.263 0.721 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.54 0.576 5.632 0.753 ;
              RECT  5.54 0.4345 5.625 0.753 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.974 0.576 5.356 0.6325 ;
              RECT  5.2995 0.548 5.356 0.6325 ;
        END
    END E
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.0725 0.576 4.26 0.799 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.012 0.4805 3.0685 0.834 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.134 0.576 0.4805 0.6325 ;
              RECT  0.134 0.569 0.4735 0.6325 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7775 0.212 0.82 0.601 ;
              RECT  0.449 0.212 0.82 0.2545 ;
              RECT  0.166 0.456 0.5935 0.4985 ;
              RECT  0.449 0.212 0.491 0.4985 ;
              RECT  0.166 0.4415 0.3075 0.4985 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.798 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.798 0.042 ;
        END
    END VSS
END SEDFFTRX2

MACRO SDFFNSRX2
    CLASS CORE ;
    SIZE 6.081 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.5755 0.643 5.6705 0.7 ;
              RECT  5.593 0.35 5.6495 0.4345 ;
              RECT  5.5755 0.378 5.632 0.7 ;
              RECT  5.54 0.4415 5.632 0.4985 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.236 0.35 5.2785 0.997 ;
              RECT  5.1335 0.6925 5.2785 0.7845 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3955 0.2965 0.4525 0.385 ;
              RECT  0.1375 0.325 0.4525 0.3815 ;
              RECT  0.325 0.2965 0.4525 0.3815 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END SE
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.4415 2.45 0.4985 ;
              RECT  2.305 0.233 2.3615 0.4985 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.4595 0.806 0.813 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5585 0.325 0.721 ;
              RECT  0.2685 0.4525 0.325 0.721 ;
        END
    END SI
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.992 0.4875 5.0485 0.841 ;
        END
    END RN
    PIN CKN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9435 0.576 1.1345 0.6325 ;
              RECT  0.9435 0.4135 1.0005 0.6325 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.081 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.081 0.042 ;
        END
    END VSS
END SDFFNSRX2

MACRO INVX8
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.05 0.509 1.1065 0.5655 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.509 0.106 0.615 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END INVX8

MACRO AOI33X1
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.6925 1.0885 0.7845 ;
              RECT  1.032 0.311 1.0745 1.0465 ;
              RECT  0.707 0.8485 1.0745 0.8905 ;
              RECT  0.562 0.311 1.0745 0.3535 ;
              RECT  0.707 0.8485 0.7495 0.933 ;
              RECT  0.562 0.2685 0.6045 0.3535 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.346 0.24 0.7 ;
        END
    END A0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.424 0.523 0.7775 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.76 0.424 0.8165 0.615 ;
              RECT  0.7495 0.5585 0.806 0.767 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.424 0.9475 0.7775 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.1625 0.3815 0.516 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.7775 ;
        END
    END B2
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END AOI33X1

MACRO OR4X4
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.269 0.7 1.3715 0.919 ;
              RECT  1.329 0.286 1.3715 0.919 ;
              RECT  1.018 0.3425 1.3715 0.385 ;
              RECT  1.308 0.286 1.3715 0.385 ;
              RECT  1.269 0.7 1.3115 0.9615 ;
              RECT  0.979 0.7 1.3715 0.742 ;
              RECT  1.018 0.286 1.0605 0.385 ;
              RECT  0.979 0.7 1.0215 0.9615 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.47 0.456 0.5265 0.6505 ;
              RECT  0.4665 0.5585 0.523 0.806 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5655 0.3955 0.795 ;
              RECT  0.339 0.456 0.3955 0.795 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.24 0.7845 ;
        END
    END D
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7105 0.4595 0.9475 0.516 ;
              RECT  0.8905 0.3425 0.9475 0.516 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END OR4X4

MACRO DFFNSRX1
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6645 0.3075 0.707 0.392 ;
              RECT  0.661 0.675 0.7035 0.951 ;
              RECT  0.629 0.3355 0.6715 0.7845 ;
              RECT  0.608 0.675 0.7035 0.7845 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.2895 0.2295 0.912 ;
              RECT  0.042 0.2895 0.2295 0.3815 ;
        END
    END QN
    PIN CKN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.285 0.3675 4.3415 0.721 ;
        END
    END CKN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.85 0.325 3.917 0.576 ;
              RECT  3.85 0.325 3.9065 0.668 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7965 0.993 3.1605 1.0355 ;
              RECT  2.7965 0.8375 2.839 1.0355 ;
              RECT  2.1955 0.8375 2.839 0.88 ;
              RECT  1.488 0.827 2.2375 0.8695 ;
              RECT  1.488 0.7105 1.5305 0.8695 ;
              RECT  1.4565 0.544 1.5025 0.767 ;
              RECT  1.4385 0.7105 1.5305 0.767 ;
              RECT  1.4175 0.544 1.5025 0.5865 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.774 0.576 0.965 0.6325 ;
              RECT  0.774 0.576 0.9475 0.795 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END DFFNSRX1

MACRO NAND3X2
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2545 0.7455 1.1065 0.788 ;
              RECT  1.064 0.2365 1.1065 0.788 ;
              RECT  1.0145 0.7105 1.1065 0.788 ;
              RECT  0.562 0.2365 1.1065 0.279 ;
              RECT  0.841 0.7455 0.8835 0.9435 ;
              RECT  0.5515 0.7455 0.5935 0.9435 ;
              RECT  0.2545 0.7455 0.304 0.9435 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3675 0.576 0.6785 0.6325 ;
              RECT  0.3675 0.576 0.5405 0.675 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.463 0.806 0.6505 ;
              RECT  0.332 0.463 0.806 0.5055 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.35 0.919 0.5195 ;
              RECT  0.219 0.35 0.919 0.392 ;
              RECT  0.1835 0.424 0.2615 0.5195 ;
              RECT  0.219 0.35 0.2615 0.5195 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END NAND3X2

MACRO ADDFHX4
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.6945 0.424 3.7755 0.516 ;
              RECT  3.355 0.707 3.737 0.7495 ;
              RECT  3.6945 0.35 3.737 0.7495 ;
              RECT  3.652 0.293 3.6945 0.392 ;
              RECT  3.645 0.707 3.6875 0.9825 ;
              RECT  3.355 0.35 3.737 0.392 ;
              RECT  3.355 0.707 3.3975 0.9825 ;
              RECT  3.355 0.293 3.3975 0.392 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.537 0.6505 0.5795 0.9155 ;
              RECT  0.1835 0.424 0.5795 0.4665 ;
              RECT  0.537 0.3675 0.5795 0.4665 ;
              RECT  0.1975 0.6505 0.5795 0.6925 ;
              RECT  0.24 0.6505 0.2825 0.9155 ;
              RECT  0.24 0.3675 0.2825 0.4665 ;
              RECT  0.1975 0.424 0.24 0.6925 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.245 0.5795 3.058 0.622 ;
              RECT  1.598 0.622 2.287 0.6645 ;
              RECT  1.598 0.5585 1.785 0.6645 ;
              RECT  1.248 0.5585 1.785 0.601 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1285 0.4415 3.171 0.5265 ;
              RECT  2.9945 0.4415 3.171 0.509 ;
              RECT  2.1315 0.4665 3.171 0.509 ;
              RECT  1.856 0.509 2.174 0.5515 ;
              RECT  1.856 0.445 1.8985 0.5515 ;
              RECT  1.0885 0.445 1.8985 0.4875 ;
              RECT  1.0885 0.445 1.131 0.53 ;
        END
    END A
    PIN CI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.955 0.3535 2.839 0.3955 ;
              RECT  1.976 0.3535 2.061 0.438 ;
              RECT  1.58 0.332 1.9975 0.3745 ;
              RECT  1.58 0.3075 1.672 0.3745 ;
        END
    END CI
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END ADDFHX4

MACRO NAND3X4
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.743 0.742 1.937 0.7845 ;
              RECT  1.895 0.286 1.937 0.7845 ;
              RECT  1.8805 0.6925 1.937 0.7845 ;
              RECT  0.6325 0.286 1.937 0.3285 ;
              RECT  1.743 0.735 1.785 0.993 ;
              RECT  0.293 0.795 1.785 0.8375 ;
              RECT  1.453 0.795 1.4955 0.993 ;
              RECT  1.163 0.795 1.2055 0.993 ;
              RECT  0.873 0.795 0.9155 0.993 ;
              RECT  0.583 0.795 0.6255 0.993 ;
              RECT  0.293 0.7175 0.3355 0.993 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.6295 0.622 1.8065 0.6645 ;
              RECT  1.764 0.5795 1.8065 0.6645 ;
              RECT  0.4525 0.682 1.672 0.7245 ;
              RECT  1.6295 0.622 1.672 0.7245 ;
              RECT  1.0425 0.6255 1.1275 0.7245 ;
              RECT  0.4525 0.6045 0.4945 0.7245 ;
              RECT  0.2155 0.6045 0.4945 0.647 ;
              RECT  0.166 0.576 0.258 0.6325 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5165 0.484 1.6935 0.5265 ;
              RECT  1.598 0.4415 1.6935 0.5265 ;
              RECT  1.598 0.424 1.6545 0.5265 ;
              RECT  1.1985 0.569 1.559 0.6115 ;
              RECT  1.5165 0.484 1.559 0.6115 ;
              RECT  1.1985 0.5125 1.2405 0.6115 ;
              RECT  0.894 0.5125 1.2405 0.555 ;
              RECT  0.5655 0.569 0.9365 0.6115 ;
              RECT  0.894 0.5125 0.9365 0.6115 ;
              RECT  0.5655 0.491 0.608 0.6115 ;
              RECT  0.364 0.491 0.608 0.5335 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3115 0.456 1.4035 0.4985 ;
              RECT  1.3115 0.3995 1.354 0.4985 ;
              RECT  0.7315 0.3995 1.354 0.4415 ;
              RECT  0.6785 0.456 0.8235 0.4985 ;
              RECT  0.7315 0.3995 0.8235 0.4985 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END NAND3X4

MACRO NOR2X8
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.061 0.6785 2.22 0.7845 ;
              RECT  2.1775 0.346 2.22 0.7845 ;
              RECT  0.226 0.346 2.22 0.3885 ;
              RECT  2.061 0.6785 2.1035 0.979 ;
              RECT  0.463 0.7035 2.22 0.7455 ;
              RECT  1.552 0.7035 1.5945 0.979 ;
              RECT  0.919 0.7035 0.9615 0.979 ;
              RECT  0.463 0.7035 0.5055 0.979 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.9125 0.5655 2.0715 0.608 ;
              RECT  0.601 0.59 1.955 0.6325 ;
              RECT  1.863 0.576 2.0715 0.608 ;
              RECT  1.4315 0.5725 1.5165 0.6325 ;
              RECT  0.997 0.5725 1.0815 0.6325 ;
              RECT  0.4875 0.5725 0.643 0.615 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.587 0.477 1.8135 0.5195 ;
              RECT  0.339 0.4595 1.6295 0.502 ;
              RECT  1.276 0.4595 1.361 0.5195 ;
              RECT  0.714 0.4595 0.799 0.5195 ;
              RECT  0.325 0.5515 0.3815 0.6505 ;
              RECT  0.339 0.4595 0.3815 0.6505 ;
              RECT  0.205 0.5515 0.3815 0.5935 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END NOR2X8

MACRO AOI32XL
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8485 0.742 0.8905 0.88 ;
              RECT  0.608 0.742 0.8905 0.7845 ;
              RECT  0.608 0.6925 0.6645 0.7845 ;
              RECT  0.622 0.3005 0.6645 0.7845 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.339 0.3955 0.629 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.1625 0.806 0.516 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.47 0.1905 0.5265 0.5055 ;
              RECT  0.4665 0.1555 0.523 0.247 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9615 0.5935 1.018 0.7915 ;
              RECT  0.8905 0.5935 1.018 0.6505 ;
              RECT  0.8905 0.509 0.9475 0.6505 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.438 0.24 0.7915 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END AOI32XL

MACRO OAI22X4
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.418 0.3145 2.5135 0.357 ;
              RECT  1.354 0.35 2.4605 0.392 ;
              RECT  2.1385 0.3145 2.2235 0.392 ;
              RECT  2.1385 0.689 2.181 0.951 ;
              RECT  0.601 0.774 2.181 0.8165 ;
              RECT  1.849 0.3145 1.9335 0.392 ;
              RECT  1.7005 0.774 1.743 0.859 ;
              RECT  1.559 0.3145 1.644 0.392 ;
              RECT  1.4385 0.774 1.5305 0.9015 ;
              RECT  1.354 0.35 1.3965 0.8165 ;
              RECT  1.085 0.7035 1.1275 0.951 ;
              RECT  0.601 0.7035 0.643 0.951 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5265 0.576 1.057 0.6325 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.725 0.576 2.2485 0.6185 ;
              RECT  1.725 0.576 1.955 0.6325 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.127 0.456 1.283 0.4985 ;
              RECT  0.873 0.4415 0.965 0.4985 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.467 0.463 2.542 0.5055 ;
              RECT  1.598 0.463 1.6545 0.6505 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END OAI22X4

MACRO OR2XL
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.5585 0.6645 0.767 ;
              RECT  0.615 0.279 0.6645 0.767 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5585 0.523 0.6785 ;
              RECT  0.3745 0.5585 0.523 0.643 ;
              RECT  0.3745 0.417 0.431 0.643 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.1905 0.615 ;
              RECT  0.134 0.417 0.1905 0.615 ;
              RECT  0.042 0.5585 0.0985 0.6785 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END OR2XL

MACRO SDFFSRHQX4
    CLASS CORE ;
    SIZE 6.081 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.905 3.6305 0.9475 ;
              RECT  2.8845 0.866 3.196 0.9085 ;
              RECT  2.319 0.951 2.927 0.993 ;
              RECT  2.8845 0.866 2.927 0.993 ;
              RECT  2.319 0.7105 2.3615 0.993 ;
              RECT  2.0435 0.7105 2.3615 0.753 ;
              RECT  2.146 0.7105 2.2375 0.767 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.883 0.4415 5.9395 0.5265 ;
              RECT  5.275 0.4415 5.9395 0.4985 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.455 0.59 5.752 0.682 ;
              RECT  5.54 0.569 5.752 0.682 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.8505 0.6115 4.9355 0.767 ;
              RECT  4.8505 0.4415 4.907 0.767 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.723 0.576 4.78 0.7565 ;
              RECT  4.55 0.576 4.78 0.6325 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.53 1.23 0.8835 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5975 0.636 0.6395 0.912 ;
              RECT  0.5975 0.371 0.6395 0.456 ;
              RECT  0.5655 0.4135 0.608 0.6785 ;
              RECT  0.3075 0.456 0.608 0.4985 ;
              RECT  0.3075 0.4415 0.3995 0.4985 ;
              RECT  0.3075 0.3815 0.35 0.912 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.081 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.081 0.042 ;
        END
    END VSS
END SDFFSRHQX4

MACRO TBUFX20
    CLASS CORE ;
    SIZE 7.071 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  6.834 0.7245 6.8765 1.0005 ;
              RECT  6.802 0.3355 6.8445 0.767 ;
              RECT  4.2565 0.7245 6.8765 0.767 ;
              RECT  6.1905 0.392 6.8445 0.4345 ;
              RECT  6.7705 0.3355 6.8445 0.4345 ;
              RECT  6.544 0.7245 6.5865 1.0005 ;
              RECT  6.4805 0.3355 6.523 0.4345 ;
              RECT  6.254 0.7245 6.2965 1.0005 ;
              RECT  6.1905 0.3355 6.233 0.4345 ;
              RECT  5.964 0.7245 6.0065 1.0005 ;
              RECT  5.9005 0.3355 5.943 0.767 ;
              RECT  5.6105 0.392 5.943 0.4345 ;
              RECT  5.6745 0.7245 5.7165 1.0005 ;
              RECT  5.6105 0.3355 5.653 0.4345 ;
              RECT  5.3845 0.7245 5.427 1.0005 ;
              RECT  5.031 0.392 5.363 0.4345 ;
              RECT  5.3205 0.3355 5.363 0.4345 ;
              RECT  5.0945 0.392 5.137 1.0005 ;
              RECT  5.031 0.3355 5.073 0.4345 ;
              RECT  4.8045 0.7245 4.847 1.0005 ;
              RECT  4.451 0.392 4.7835 0.4345 ;
              RECT  4.741 0.3355 4.7835 0.4345 ;
              RECT  4.5145 0.392 4.557 1.0005 ;
              RECT  4.451 0.3355 4.4935 0.4345 ;
              RECT  4.2565 0.424 4.3415 0.516 ;
              RECT  4.2565 0.424 4.299 0.7845 ;
              RECT  4.2245 0.742 4.267 1.0005 ;
              RECT  4.161 0.424 4.3415 0.4665 ;
              RECT  4.161 0.3355 4.2035 0.4665 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.018 0.576 1.4565 0.6185 ;
              RECT  1.414 0.516 1.4565 0.6185 ;
              RECT  1.156 0.576 1.248 0.6325 ;
              RECT  1.018 0.516 1.0605 0.6185 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.16 0.484 3.9275 0.5265 ;
              RECT  2.16 0.392 2.2025 0.5265 ;
              RECT  2.135 0.2435 2.1775 0.4345 ;
              RECT  1.8665 0.2435 2.1775 0.286 ;
              RECT  1.64 0.392 1.909 0.4345 ;
              RECT  1.8665 0.2435 1.909 0.4345 ;
              RECT  1.7075 0.392 1.75 0.5335 ;
              RECT  1.64 0.212 1.6825 0.4345 ;
              RECT  1.361 0.212 1.6825 0.2545 ;
              RECT  1.1345 0.392 1.4035 0.4345 ;
              RECT  1.361 0.212 1.4035 0.4345 ;
              RECT  1.209 0.392 1.2515 0.5055 ;
              RECT  1.1345 0.212 1.177 0.4345 ;
              RECT  0.7175 0.212 1.177 0.2545 ;
              RECT  0.491 0.41 0.76 0.4525 ;
              RECT  0.7175 0.212 0.76 0.4525 ;
              RECT  0.6645 0.41 0.707 0.509 ;
              RECT  0.5515 0.41 0.5935 0.509 ;
              RECT  0.491 0.212 0.5335 0.4525 ;
              RECT  0.1975 0.212 0.5335 0.2545 ;
              RECT  0.1975 0.212 0.24 0.484 ;
              RECT  0.0245 0.4415 0.1975 0.4985 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 7.071 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 7.071 0.042 ;
        END
    END VSS
END TBUFX20

MACRO INVX16
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.0645 0.4985 2.121 0.5655 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.509 0.106 0.615 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END INVX16

MACRO ADDHX4
    CLASS CORE ;
    SIZE 2.9695 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.57 0.576 2.6125 0.721 ;
              RECT  2.1705 0.403 2.588 0.445 ;
              RECT  2.1775 0.576 2.6125 0.6185 ;
              RECT  2.305 0.5585 2.3615 0.6505 ;
              RECT  2.319 0.403 2.3615 0.6505 ;
              RECT  2.1775 0.576 2.22 0.8835 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.905 0.7565 1.0605 0.799 ;
              RECT  0.5655 0.41 1.0605 0.4525 ;
              RECT  1.018 0.3605 1.0605 0.4525 ;
              RECT  0.905 0.41 0.9475 0.799 ;
              RECT  0.643 0.6715 0.9475 0.714 ;
              RECT  0.8905 0.41 0.9475 0.714 ;
              RECT  0.5655 0.3675 0.608 0.4525 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.291 0.7915 2.786 0.834 ;
              RECT  2.7435 0.523 2.786 0.834 ;
              RECT  2.291 0.7915 2.333 0.997 ;
              RECT  1.8985 0.9545 2.333 0.997 ;
              RECT  1.3575 0.972 1.941 1.0145 ;
              RECT  1.347 0.5515 1.4315 0.5935 ;
              RECT  1.3575 0.5515 1.4 1.0145 ;
              RECT  0.5795 0.8695 1.4 0.912 ;
              RECT  0.5795 0.806 0.622 0.912 ;
              RECT  0.0985 0.806 0.622 0.8485 ;
              RECT  0.0985 0.537 0.141 0.8485 ;
              RECT  0.042 0.5585 0.141 0.6505 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.131 0.438 1.3115 0.4805 ;
              RECT  1.131 0.247 1.1735 0.4805 ;
              RECT  0.905 0.247 1.1735 0.2895 ;
              RECT  0.4525 0.2545 0.9475 0.2965 ;
              RECT  0.325 0.424 0.4945 0.4665 ;
              RECT  0.4525 0.2545 0.4945 0.4665 ;
              RECT  0.325 0.424 0.3815 0.5655 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.9695 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.9695 0.042 ;
        END
    END VSS
END ADDHX4

MACRO SDFFSHQX8
    CLASS CORE ;
    SIZE 5.6565 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.774 0.6575 1.1875 0.7 ;
              RECT  1.1455 0.3815 1.1875 0.7 ;
              RECT  1.064 0.6575 1.1065 0.742 ;
              RECT  0.774 0.3815 0.8165 0.951 ;
              RECT  0.7495 0.424 0.8165 0.516 ;
              RECT  0.194 0.424 0.8165 0.4665 ;
              RECT  0.484 0.3815 0.5265 0.951 ;
              RECT  0.194 0.3815 0.2365 0.951 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.5575 0.5585 5.614 0.6505 ;
              RECT  4.9815 0.516 5.6 0.5585 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.176 0.668 5.487 0.767 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4085 0.5725 4.6735 0.629 ;
              RECT  4.4085 0.4945 4.5005 0.6395 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.267 0.7105 4.43 0.767 ;
              RECT  4.267 0.5335 4.338 0.767 ;
              RECT  4.253 0.5335 4.338 0.59 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.669 0.6715 2.786 0.714 ;
              RECT  2.485 0.8625 2.7115 0.905 ;
              RECT  2.669 0.6715 2.7115 0.905 ;
              RECT  1.771 0.912 2.5275 0.9545 ;
              RECT  2.485 0.8625 2.5275 0.9545 ;
              RECT  1.771 0.6575 1.8205 0.742 ;
              RECT  1.771 0.6575 1.8135 0.9545 ;
              RECT  1.7215 0.7105 1.8135 0.767 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.6565 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.6565 0.042 ;
        END
    END VSS
END SDFFSHQX8

MACRO DFFRHQX2
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3745 0.24 0.9225 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.576 1.248 0.6325 ;
              RECT  1.05 0.7245 1.2125 0.788 ;
              RECT  1.156 0.576 1.2125 0.788 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.424 0.7105 0.59 0.767 ;
              RECT  0.424 0.523 0.5405 0.767 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8955 0.364 2.952 0.6255 ;
              RECT  2.8035 0.364 2.952 0.4985 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END DFFRHQX2

MACRO DFFNSRX4
    CLASS CORE ;
    SIZE 5.515 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.663 0.357 5.0805 0.3995 ;
              RECT  4.8715 0.608 4.914 0.94 ;
              RECT  4.426 0.608 4.914 0.6505 ;
              RECT  4.663 0.357 4.7055 0.6505 ;
              RECT  4.582 0.608 4.624 0.94 ;
              RECT  4.426 0.5585 4.483 0.6505 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.9985 0.357 4.4155 0.3995 ;
              RECT  4.292 0.7105 4.3345 0.94 ;
              RECT  3.9845 0.7105 4.3345 0.753 ;
              RECT  4.041 0.357 4.0835 0.753 ;
              RECT  3.9845 0.7105 4.076 0.767 ;
              RECT  3.9845 0.7105 4.0265 0.94 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.04 0.445 2.206 0.502 ;
              RECT  1.983 0.576 2.0965 0.6325 ;
              RECT  2.04 0.445 2.0965 0.6325 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.58 0.47 1.9055 0.5265 ;
              RECT  1.58 0.4415 1.672 0.5265 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.537 0.3815 0.8905 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.537 0.24 0.8905 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.515 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.515 0.042 ;
        END
    END VSS
END DFFNSRX4

MACRO TLATNSRX4
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.3695 0.608 4.412 0.9295 ;
              RECT  4.1115 0.608 4.412 0.6505 ;
              RECT  4.023 0.438 4.3555 0.4805 ;
              RECT  4.313 0.3815 4.3555 0.4805 ;
              RECT  4.1115 0.438 4.2 0.6505 ;
              RECT  4.1115 0.438 4.154 0.7035 ;
              RECT  4.08 0.661 4.122 0.9295 ;
              RECT  4.023 0.3815 4.0655 0.4805 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.164 0.654 3.2065 0.9295 ;
              RECT  2.8635 0.438 3.196 0.4805 ;
              RECT  3.1535 0.3815 3.196 0.4805 ;
              RECT  2.8705 0.654 3.2065 0.6965 ;
              RECT  2.8845 0.438 2.927 0.7845 ;
              RECT  2.8705 0.654 2.9165 0.9295 ;
              RECT  2.8635 0.3815 2.906 0.4805 ;
        END
    END QN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.57 0.555 2.6795 0.5975 ;
              RECT  2.57 0.555 2.662 0.6325 ;
              RECT  2.2235 0.6185 2.6125 0.661 ;
              RECT  2.2235 0.562 2.266 0.661 ;
              RECT  2.181 0.562 2.266 0.6045 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.491 1.23 0.8445 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0355 0.212 2.075 0.2545 ;
              RECT  1.0355 0.152 1.078 0.2545 ;
              RECT  0.5865 0.152 1.078 0.194 ;
              RECT  0.449 0.576 0.629 0.6325 ;
              RECT  0.5865 0.152 0.629 0.6325 ;
              RECT  0.311 0.576 0.629 0.6185 ;
        END
    END RN
    PIN GN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.4945 0.24 0.8485 ;
        END
    END GN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END TLATNSRX4

MACRO ADDFHX2
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.136 0.424 3.21 0.516 ;
              RECT  3.136 0.3815 3.178 0.767 ;
              RECT  3.104 0.7245 3.1465 0.9825 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.3815 0.24 0.912 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.075 0.5795 2.807 0.622 ;
              RECT  1.2975 0.6395 2.1175 0.682 ;
              RECT  2.075 0.5795 2.1175 0.682 ;
              RECT  1.2975 0.6395 1.389 0.767 ;
              RECT  0.965 0.6045 1.3395 0.647 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8775 0.4665 2.92 0.5515 ;
              RECT  1.962 0.4665 2.92 0.509 ;
              RECT  2.7115 0.4415 2.8035 0.509 ;
              RECT  1.7005 0.5265 2.0045 0.569 ;
              RECT  1.962 0.4665 2.0045 0.569 ;
              RECT  0.8695 0.491 1.743 0.5335 ;
              RECT  0.8095 0.4945 0.894 0.537 ;
        END
    END A
    PIN CI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.831 0.3535 2.595 0.3955 ;
              RECT  1.831 0.3535 1.8735 0.456 ;
              RECT  1.2975 0.371 1.8735 0.4135 ;
              RECT  1.2975 0.3075 1.389 0.4135 ;
        END
    END CI
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END ADDFHX2

MACRO NOR4BBXL
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.5585 0.9475 0.6505 ;
              RECT  0.523 0.9545 0.933 0.997 ;
              RECT  0.8905 0.18 0.933 0.997 ;
              RECT  0.5865 0.318 0.933 0.3605 ;
              RECT  0.5865 0.18 0.629 0.3605 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4805 0.544 0.537 0.813 ;
              RECT  0.4665 0.6925 0.523 0.8835 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.6925 0.767 0.7915 ;
              RECT  0.7105 0.544 0.767 0.7915 ;
              RECT  0.608 0.6925 0.6645 0.795 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.576 1.248 0.6325 ;
              RECT  1.078 0.76 1.2125 0.8165 ;
              RECT  1.156 0.576 1.2125 0.8165 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.021 0.484 0.2825 0.6325 ;
        END
    END BN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END NOR4BBXL

MACRO NOR2X6
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.41 0.7245 1.6825 0.767 ;
              RECT  1.64 0.35 1.6825 0.767 ;
              RECT  1.598 0.6925 1.6545 0.7845 ;
              RECT  0.194 0.35 1.6825 0.392 ;
              RECT  1.354 0.7245 1.3965 0.9435 ;
              RECT  1.354 0.3075 1.3965 0.392 ;
              RECT  1.064 0.3075 1.1065 0.392 ;
              RECT  0.866 0.7245 0.9085 0.9435 ;
              RECT  0.774 0.3075 0.8165 0.392 ;
              RECT  0.484 0.3075 0.5265 0.392 ;
              RECT  0.41 0.7245 0.4525 0.9435 ;
              RECT  0.194 0.3075 0.2365 0.392 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2975 0.576 1.4565 0.6325 ;
              RECT  0.548 0.6045 1.3325 0.647 ;
              RECT  0.8165 0.576 0.9015 0.647 ;
              RECT  0.4345 0.576 0.59 0.6185 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.527 0.463 1.5695 0.622 ;
              RECT  0.1975 0.463 1.5695 0.5055 ;
              RECT  1.096 0.463 1.1805 0.5335 ;
              RECT  0.661 0.463 0.7455 0.5335 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
              RECT  0.1975 0.463 0.24 0.6505 ;
              RECT  0.152 0.5585 0.24 0.601 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END NOR2X6

MACRO CLKBUFX8
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.997 0.3885 1.092 0.431 ;
              RECT  1.0285 0.6575 1.071 0.972 ;
              RECT  0.159 0.3995 1.0285 0.4415 ;
              RECT  0.159 0.6575 1.071 0.7 ;
              RECT  0.7175 0.3885 0.8025 0.4415 ;
              RECT  0.7385 0.6575 0.781 0.972 ;
              RECT  0.4275 0.3885 0.5125 0.4415 ;
              RECT  0.449 0.6575 0.491 0.972 ;
              RECT  0.1835 0.3995 0.24 0.516 ;
              RECT  0.1835 0.3995 0.226 0.7 ;
              RECT  0.159 0.6575 0.2015 0.972 ;
              RECT  0.159 0.357 0.2015 0.4415 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4565 0.424 1.513 0.7775 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END CLKBUFX8

MACRO NOR2BX4
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0245 0.346 1.1065 0.3885 ;
              RECT  1.064 0.304 1.1065 0.3885 ;
              RECT  0.8165 0.7035 0.859 0.9615 ;
              RECT  0.774 0.304 0.8165 0.3885 ;
              RECT  0.0245 0.7035 0.859 0.7455 ;
              RECT  0.484 0.304 0.5265 0.3885 ;
              RECT  0.378 0.7035 0.4205 0.9615 ;
              RECT  0.194 0.304 0.2365 0.3885 ;
              RECT  0.0245 0.576 0.1165 0.6325 ;
              RECT  0.0245 0.346 0.067 0.7455 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.41 0.576 0.8835 0.6325 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.6925 1.2515 0.7495 ;
              RECT  1.195 0.5725 1.2515 0.7495 ;
              RECT  1.032 0.6925 1.0885 0.7845 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END NOR2BX4

MACRO TLATNSRX1
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.622 0.2895 0.6645 0.94 ;
              RECT  0.608 0.2895 0.6645 0.3815 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.159 0.3815 0.2155 0.912 ;
              RECT  0.042 0.424 0.2155 0.516 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8705 0.6925 3.0015 0.7495 ;
              RECT  2.945 0.555 3.0015 0.7495 ;
              RECT  2.8705 0.6925 2.927 0.834 ;
        END
    END GN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.6195 0.5975 2.8 0.6395 ;
              RECT  2.57 0.576 2.662 0.6325 ;
              RECT  2.6195 0.212 2.662 0.6395 ;
              RECT  1.269 0.212 2.662 0.2545 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.022 0.438 2.0785 0.6505 ;
              RECT  1.994 0.5655 2.0505 0.7635 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8485 0.5725 0.9475 0.629 ;
              RECT  0.7495 0.6925 0.905 0.7845 ;
              RECT  0.8485 0.5725 0.905 0.7845 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END TLATNSRX1

MACRO AOI2BB1XL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2225 0.2015 0.318 0.2435 ;
              RECT  0.0565 0.318 0.265 0.3605 ;
              RECT  0.2225 0.2015 0.265 0.3605 ;
              RECT  0.18 0.608 0.2225 0.979 ;
              RECT  0.042 0.608 0.2225 0.6505 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
              RECT  0.0565 0.318 0.0985 0.6505 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.332 0.544 0.3885 0.7495 ;
              RECT  0.325 0.6925 0.3815 0.8905 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4595 0.6925 0.523 0.8905 ;
              RECT  0.4595 0.544 0.516 0.8905 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.707 0.318 0.806 0.6715 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END AOI2BB1XL

MACRO NOR3X8
    CLASS CORE ;
    SIZE 3.6765 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4715 0.7105 3.652 0.767 ;
              RECT  0.24 0.194 3.6485 0.2365 ;
              RECT  3.4715 0.636 3.5955 0.767 ;
              RECT  3.553 0.194 3.5955 0.767 ;
              RECT  3.4715 0.636 3.514 0.951 ;
              RECT  0.707 0.7705 3.514 0.813 ;
              RECT  2.662 0.7705 2.7045 0.8555 ;
              RECT  1.5905 0.7705 1.633 0.8555 ;
              RECT  0.707 0.7705 0.7495 0.8555 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9625 0.544 3.0475 0.5865 ;
              RECT  0.364 0.6575 3.005 0.7 ;
              RECT  2.9625 0.544 3.005 0.7 ;
              RECT  2.001 0.544 2.0855 0.5865 ;
              RECT  2.001 0.544 2.0435 0.7 ;
              RECT  1.191 0.544 1.2335 0.7 ;
              RECT  1.149 0.544 1.2335 0.5865 ;
              RECT  0.364 0.59 0.4065 0.7 ;
              RECT  0.166 0.59 0.4065 0.6325 ;
              RECT  0.166 0.576 0.2615 0.6325 ;
              RECT  0.219 0.516 0.2615 0.6325 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.277 0.4415 3.369 0.4985 ;
              RECT  3.118 0.4415 3.369 0.484 ;
              RECT  2.8495 0.431 3.1605 0.4735 ;
              RECT  2.768 0.438 2.892 0.4805 ;
              RECT  2.4995 0.544 2.8105 0.5865 ;
              RECT  2.768 0.438 2.8105 0.5865 ;
              RECT  2.4995 0.438 2.542 0.5865 ;
              RECT  2.287 0.438 2.542 0.4805 ;
              RECT  1.8525 0.431 2.3295 0.4735 ;
              RECT  1.81 0.438 1.895 0.4805 ;
              RECT  1.5025 0.544 1.8525 0.5865 ;
              RECT  1.81 0.438 1.8525 0.5865 ;
              RECT  1.5025 0.431 1.545 0.5865 ;
              RECT  0.894 0.431 1.545 0.4735 ;
              RECT  1.3505 0.431 1.393 0.516 ;
              RECT  0.852 0.438 0.9365 0.4805 ;
              RECT  0.477 0.544 0.894 0.5865 ;
              RECT  0.852 0.438 0.894 0.5865 ;
              RECT  0.477 0.477 0.5195 0.5865 ;
              RECT  0.332 0.477 0.5195 0.5195 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.44 0.3075 3.4825 0.5125 ;
              RECT  0.59 0.3075 3.4825 0.35 ;
              RECT  2.6125 0.431 2.6975 0.4735 ;
              RECT  2.6125 0.3075 2.655 0.4735 ;
              RECT  1.6155 0.431 1.7005 0.4735 ;
              RECT  1.658 0.3075 1.7005 0.4735 ;
              RECT  0.59 0.3075 0.7565 0.4735 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.6765 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.6765 0.042 ;
        END
    END VSS
END NOR3X8

MACRO ADDHX2
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.643 1.704 0.7 ;
              RECT  1.598 0.371 1.6545 0.7 ;
              RECT  1.5625 0.371 1.6545 0.4275 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6115 0.7315 0.806 0.788 ;
              RECT  0.7495 0.392 0.806 0.788 ;
              RECT  0.544 0.392 0.806 0.449 ;
        END
    END CO
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.919 0.905 0.9615 0.9895 ;
              RECT  0.601 0.905 0.9615 0.9475 ;
              RECT  0.601 0.859 0.643 0.9475 ;
              RECT  0.4985 0.859 0.643 0.9015 ;
              RECT  0.4985 0.6325 0.5405 0.9015 ;
              RECT  0.4345 0.6325 0.5405 0.767 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.258 1.969 0.3005 ;
              RECT  1.209 0.1625 1.294 0.3005 ;
              RECT  1.032 0.258 1.0745 0.6785 ;
              RECT  0.1835 0.424 0.24 0.5865 ;
              RECT  0.1835 0.258 0.226 0.5865 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END ADDHX2

MACRO SDFFSHQX2
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2965 0.3605 0.3535 0.912 ;
              RECT  0.166 0.4415 0.3535 0.4985 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.426 0.424 4.483 0.516 ;
              RECT  3.9065 0.449 4.483 0.5055 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.062 0.576 4.3555 0.6325 ;
              RECT  4.062 0.576 4.1185 0.6925 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4365 0.4415 3.521 0.5585 ;
              RECT  3.2275 0.4415 3.521 0.4985 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.224 0.629 3.4965 0.6855 ;
              RECT  3.224 0.629 3.369 0.767 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.757 0.682 1.842 0.7245 ;
              RECT  0.781 0.8375 1.7995 0.88 ;
              RECT  1.757 0.682 1.7995 0.88 ;
              RECT  0.781 0.576 0.8235 0.88 ;
              RECT  0.7315 0.576 0.8235 0.6325 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END SDFFSHQX2

MACRO OAI32X4
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.026 0.3425 3.1215 0.385 ;
              RECT  2.167 0.378 3.0685 0.4205 ;
              RECT  2.747 0.3425 2.8315 0.4205 ;
              RECT  2.7365 0.8165 2.7785 0.9015 ;
              RECT  0.6395 0.8165 2.7785 0.859 ;
              RECT  2.457 0.3425 2.542 0.4205 ;
              RECT  2.298 0.8165 2.3405 0.9015 ;
              RECT  2.167 0.3425 2.252 0.4205 ;
              RECT  2.0185 0.484 2.2095 0.5265 ;
              RECT  2.167 0.3425 2.2095 0.5265 ;
              RECT  2.0185 0.484 2.061 0.859 ;
              RECT  1.7215 0.8165 1.8135 0.9015 ;
              RECT  1.5235 0.8165 1.566 0.9015 ;
              RECT  0.6395 0.8165 0.682 0.9015 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.226 0.7035 1.948 0.7455 ;
              RECT  1.9055 0.6045 1.948 0.7455 ;
              RECT  1.0075 0.6255 1.092 0.7455 ;
              RECT  0.226 0.576 0.2685 0.7455 ;
              RECT  0.166 0.576 0.2685 0.6325 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9095 0.6045 3.0685 0.6505 ;
              RECT  3.012 0.5585 3.0685 0.6505 ;
              RECT  2.1315 0.7035 2.952 0.7455 ;
              RECT  2.9095 0.6045 2.952 0.7455 ;
              RECT  2.542 0.6255 2.6265 0.7455 ;
              RECT  2.1315 0.5975 2.174 0.7455 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2725 0.59 1.8275 0.6325 ;
              RECT  1.2725 0.5125 1.315 0.6325 ;
              RECT  0.894 0.5125 1.315 0.555 ;
              RECT  0.339 0.576 0.9365 0.6185 ;
              RECT  0.894 0.5125 0.9365 0.6185 ;
              RECT  0.449 0.576 0.5405 0.6325 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7115 0.548 2.8315 0.6325 ;
              RECT  2.3295 0.5125 2.754 0.555 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4245 0.3995 1.467 0.5195 ;
              RECT  0.781 0.3995 1.467 0.4415 ;
              RECT  0.647 0.456 0.8235 0.4985 ;
              RECT  0.7315 0.4415 0.8235 0.4985 ;
        END
    END A2
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END OAI32X4

MACRO NAND4BXL
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3955 0.8165 0.608 0.859 ;
              RECT  0.3955 0.7495 0.438 0.859 ;
              RECT  0.0565 0.7495 0.438 0.7915 ;
              RECT  0.24 0.7495 0.325 0.859 ;
              RECT  0.042 0.212 0.194 0.2545 ;
              RECT  0.152 0.1695 0.194 0.2545 ;
              RECT  0.0565 0.212 0.0985 0.7915 ;
              RECT  0.042 0.212 0.0985 0.3815 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7315 0.548 0.8235 0.6325 ;
              RECT  0.7315 0.548 0.788 0.866 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.1625 0.523 0.516 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.424 0.3955 0.516 ;
              RECT  0.325 0.1765 0.3815 0.516 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.325 0.24 0.6785 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END NAND4BXL

MACRO TLATNCAX16
    CLASS CORE ;
    SIZE 5.091 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1775 0.403 2.273 0.445 ;
              RECT  0.41 0.714 2.234 0.7565 ;
              RECT  1.9195 0.4135 2.2095 0.456 ;
              RECT  1.9195 0.371 1.962 0.7565 ;
              RECT  1.598 0.403 1.6935 0.445 ;
              RECT  1.598 0.5585 1.6545 0.7565 ;
              RECT  1.598 0.403 1.64 0.7565 ;
              RECT  1.3185 0.403 1.4035 0.445 ;
              RECT  1.3185 0.403 1.3645 0.7565 ;
              RECT  1.0285 0.403 1.1135 0.445 ;
              RECT  1.0285 0.403 1.071 0.7565 ;
              RECT  0.7385 0.403 0.8235 0.445 ;
              RECT  0.7385 0.403 0.781 0.7565 ;
              RECT  0.47 0.3815 0.5125 0.7565 ;
        END
    END ECK
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.709 0.4735 4.794 0.714 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.233 0.4595 0.3815 0.516 ;
              RECT  0.325 0.424 0.3815 0.516 ;
              RECT  0.233 0.4595 0.2895 0.6855 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.091 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.091 0.042 ;
        END
    END VSS
END TLATNCAX16

MACRO FILL1
    CLASS CORE ;
    SIZE 0.141 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.141 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.141 0.042 ;
        END
    END VSS
END FILL1

MACRO DFFSHQX2
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3815 0.24 0.912 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.277 0.502 3.3725 0.6965 ;
              RECT  3.157 0.502 3.3725 0.5585 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9945 0.502 3.0865 0.742 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.036 0.456 2.0785 0.5795 ;
              RECT  1.8805 0.456 2.0785 0.4985 ;
              RECT  1.8805 0.247 1.923 0.4985 ;
              RECT  1.032 0.247 1.923 0.2895 ;
              RECT  1.032 0.424 1.0885 0.516 ;
              RECT  0.827 0.608 1.0745 0.6505 ;
              RECT  1.032 0.247 1.0745 0.6505 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END DFFSHQX2

MACRO TBUFX3
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.442 0.339 1.7745 0.3815 ;
              RECT  1.732 0.2825 1.7745 0.3815 ;
              RECT  1.725 0.636 1.7675 0.912 ;
              RECT  1.598 0.636 1.7675 0.6785 ;
              RECT  1.598 0.5585 1.6545 0.6785 ;
              RECT  1.393 0.7845 1.64 0.827 ;
              RECT  1.598 0.339 1.64 0.827 ;
              RECT  1.442 0.2825 1.4845 0.3815 ;
              RECT  1.393 0.7845 1.435 0.8695 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.184 0.1905 1.2265 0.4875 ;
              RECT  0.59 0.1905 1.2265 0.233 ;
              RECT  0.59 0.576 0.682 0.6325 ;
              RECT  0.59 0.1905 0.6325 0.6325 ;
              RECT  0.311 0.5865 0.682 0.629 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.4595 0.5195 0.516 ;
              RECT  0.1835 0.424 0.24 0.544 ;
        END
    END OE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END TBUFX3

MACRO NOR2BX2
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6575 0.325 0.742 0.3675 ;
              RECT  0.0565 0.339 0.6925 0.3815 ;
              RECT  0.4945 0.608 0.537 0.9615 ;
              RECT  0.042 0.608 0.537 0.6505 ;
              RECT  0.346 0.325 0.431 0.3815 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
              RECT  0.0565 0.339 0.0985 0.6505 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6925 0.919 0.7495 ;
              RECT  0.8625 0.5655 0.919 0.7495 ;
              RECT  0.7495 0.6925 0.806 0.806 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.5655 0.6645 0.919 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END NOR2BX2

MACRO AOI21X4
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7465 0.675 1.7885 0.76 ;
              RECT  1.4565 0.675 1.7885 0.7175 ;
              RECT  1.658 0.3145 1.743 0.357 ;
              RECT  0.6045 0.3285 1.6935 0.371 ;
              RECT  1.4565 0.576 1.5305 0.76 ;
              RECT  1.336 0.576 1.5305 0.6325 ;
              RECT  1.3785 0.286 1.421 0.371 ;
              RECT  1.336 0.3285 1.3785 0.6325 ;
              RECT  0.993 0.3145 1.078 0.371 ;
              RECT  0.555 0.3145 0.6395 0.357 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5055 0.576 1.025 0.6325 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.463 1.23 0.6505 ;
              RECT  0.3815 0.463 1.23 0.5055 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4495 0.449 1.796 0.5055 ;
              RECT  1.58 0.4415 1.672 0.5055 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END AOI21X4

MACRO OR2X6
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.919 0.424 1.541 0.4665 ;
              RECT  1.499 0.247 1.541 0.4665 ;
              RECT  1.446 0.6785 1.488 1.011 ;
              RECT  0.866 0.6785 1.488 0.721 ;
              RECT  1.315 0.424 1.3715 0.516 ;
              RECT  1.315 0.424 1.3575 0.721 ;
              RECT  1.209 0.247 1.2515 0.4665 ;
              RECT  1.156 0.6785 1.1985 1.011 ;
              RECT  0.919 0.247 0.9615 0.4665 ;
              RECT  0.866 0.6785 0.9085 1.011 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.643 0.47 0.7 ;
              RECT  0.325 0.643 0.3815 0.919 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.516 0.682 0.5725 ;
              RECT  0.1835 0.544 0.2545 0.601 ;
              RECT  0.1835 0.544 0.24 0.6505 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END OR2X6

MACRO OAI22X2
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0745 0.3145 1.17 0.357 ;
              RECT  0.7775 0.35 1.117 0.392 ;
              RECT  0.993 0.7245 1.0355 0.958 ;
              RECT  0.4525 0.7245 1.0355 0.767 ;
              RECT  0.7775 0.3145 0.88 0.392 ;
              RECT  0.661 0.4415 0.82 0.484 ;
              RECT  0.7775 0.3145 0.82 0.484 ;
              RECT  0.59 0.7105 0.7035 0.767 ;
              RECT  0.661 0.4415 0.7035 0.767 ;
              RECT  0.4525 0.7245 0.4945 0.958 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.569 0.463 0.6255 ;
              RECT  0.1835 0.569 0.24 0.7845 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.59 1.23 0.788 ;
              RECT  1.018 0.59 1.23 0.647 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5335 0.4415 0.59 0.5265 ;
              RECT  0.141 0.4415 0.59 0.4985 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.463 1.223 0.5195 ;
              RECT  0.8905 0.463 0.9475 0.6505 ;
              RECT  0.774 0.555 0.9475 0.6115 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END OAI22X2

MACRO TBUFX1
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.322 0.643 1.389 0.919 ;
              RECT  1.347 0.3075 1.389 0.919 ;
              RECT  1.2265 0.3075 1.389 0.392 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8695 0.2015 1.011 0.2435 ;
              RECT  0.509 0.219 0.912 0.2615 ;
              RECT  0.304 0.7105 0.622 0.753 ;
              RECT  0.5795 0.47 0.622 0.753 ;
              RECT  0.509 0.47 0.622 0.5125 ;
              RECT  0.509 0.219 0.5515 0.5125 ;
              RECT  0.449 0.7105 0.5405 0.767 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1765 0.583 0.509 0.6395 ;
              RECT  0.325 0.424 0.3815 0.6395 ;
              RECT  0.1765 0.583 0.233 0.668 ;
        END
    END OE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END TBUFX1

MACRO SDFFX4
    CLASS CORE ;
    SIZE 4.9495 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.009 0.346 4.426 0.3885 ;
              RECT  4.306 0.636 4.3485 0.912 ;
              RECT  4.002 0.636 4.3485 0.6785 ;
              RECT  4.002 0.5585 4.0585 0.912 ;
              RECT  4.009 0.346 4.0585 0.912 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.726 0.636 3.7685 0.912 ;
              RECT  3.3445 0.346 3.7615 0.3885 ;
              RECT  3.4365 0.636 3.7685 0.6785 ;
              RECT  3.4505 0.346 3.493 0.6785 ;
              RECT  3.4365 0.5585 3.4785 0.912 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.4525 1.248 0.6325 ;
              RECT  1.018 0.4525 1.248 0.509 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.2685 0.9475 0.622 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.4665 0.7845 ;
              RECT  0.41 0.5585 0.4665 0.7845 ;
              RECT  0.325 0.6925 0.3815 0.827 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.537 0.424 0.5935 0.6785 ;
              RECT  0.1835 0.424 0.5935 0.4875 ;
              RECT  0.279 0.403 0.3355 0.4875 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.9495 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.9495 0.042 ;
        END
    END VSS
END SDFFX4

MACRO INVX12
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4845 0.4985 1.541 0.5655 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.509 0.106 0.615 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END INVX12

MACRO DFFRHQX8
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.55 0.449 4.642 0.767 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.686 0.2435 1.7285 0.5725 ;
              RECT  1.2335 0.2435 1.7285 0.286 ;
              RECT  1.1735 0.424 1.276 0.562 ;
              RECT  1.2335 0.2435 1.276 0.562 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.122 0.332 4.366 0.4345 ;
              RECT  4.122 0.332 4.2175 0.4985 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.887 0.403 0.9895 0.445 ;
              RECT  0.919 0.636 0.9615 0.951 ;
              RECT  0.887 0.403 0.9295 0.6785 ;
              RECT  0.629 0.523 0.9295 0.5655 ;
              RECT  0.636 0.3815 0.6785 0.5655 ;
              RECT  0.629 0.4735 0.6715 0.951 ;
              RECT  0.042 0.4735 0.6785 0.516 ;
              RECT  0.346 0.3815 0.3885 0.516 ;
              RECT  0.339 0.4735 0.3815 0.951 ;
              RECT  0.042 0.3815 0.0985 0.516 ;
              RECT  0.042 0.3815 0.0915 0.951 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END DFFRHQX8

MACRO NOR2X4
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.523 0.7035 1.389 0.7455 ;
              RECT  1.347 0.35 1.389 0.7455 ;
              RECT  1.2975 0.576 1.389 0.6325 ;
              RECT  0.3075 0.35 1.389 0.392 ;
              RECT  1.177 0.3075 1.2195 0.392 ;
              RECT  0.993 0.7035 1.0355 0.951 ;
              RECT  0.887 0.3075 0.9295 0.392 ;
              RECT  0.5975 0.3075 0.6395 0.392 ;
              RECT  0.523 0.7035 0.5655 0.951 ;
              RECT  0.3075 0.3075 0.35 0.392 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.53 0.576 1.004 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.258 0.463 1.269 0.5055 ;
              RECT  0.325 0.463 0.3815 0.6505 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END NOR2X4

MACRO OR3X8
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.075 0.403 2.16 0.445 ;
              RECT  1.2585 0.4135 2.107 0.456 ;
              RECT  2.0255 0.6395 2.068 0.951 ;
              RECT  1.156 0.6395 2.068 0.682 ;
              RECT  1.8805 0.4135 1.937 0.516 ;
              RECT  1.8805 0.4135 1.923 0.682 ;
              RECT  1.8065 0.371 1.849 0.456 ;
              RECT  1.7355 0.6395 1.778 0.951 ;
              RECT  1.4955 0.403 1.58 0.456 ;
              RECT  1.446 0.6395 1.488 0.951 ;
              RECT  1.2055 0.403 1.29 0.445 ;
              RECT  1.156 0.6395 1.1985 0.951 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.583 0.675 0.6395 ;
              RECT  0.4665 0.583 0.523 0.7845 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.47 0.8445 0.555 ;
              RECT  0.7495 0.47 0.806 0.6505 ;
              RECT  0.3745 0.47 0.8445 0.5125 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.919 0.357 0.9615 0.5335 ;
              RECT  0.2085 0.357 0.9615 0.3995 ;
              RECT  0.1835 0.3675 0.24 0.516 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END OR3X8

MACRO BUFX2
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.247 0.6115 0.2895 0.933 ;
              RECT  0.247 0.35 0.2895 0.4345 ;
              RECT  0.2155 0.392 0.258 0.654 ;
              RECT  0.1835 0.424 0.258 0.516 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3605 0.7105 0.5405 0.767 ;
              RECT  0.484 0.537 0.5405 0.767 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END BUFX2

MACRO NOR4X8
    CLASS CORE ;
    SIZE 4.384 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.154 0.576 4.1965 0.951 ;
              RECT  3.7475 0.576 4.1965 0.6185 ;
              RECT  0.2365 0.332 4.0515 0.3745 ;
              RECT  4.009 0.2895 4.0515 0.3745 ;
              RECT  3.882 0.332 3.924 0.6185 ;
              RECT  3.7475 0.576 3.917 0.6505 ;
              RECT  3.8605 0.5585 3.9065 0.8375 ;
              RECT  3.2845 0.7035 3.9065 0.7455 ;
              RECT  3.7475 0.576 3.9065 0.7455 ;
              RECT  3.698 0.3215 3.783 0.3745 ;
              RECT  3.574 0.7035 3.6165 0.8375 ;
              RECT  3.408 0.3215 3.493 0.3745 ;
              RECT  3.2845 0.7035 3.3265 0.8375 ;
              RECT  3.118 0.3215 3.203 0.3745 ;
              RECT  2.828 0.3215 2.913 0.3745 ;
              RECT  2.5385 0.3215 2.623 0.3745 ;
              RECT  2.2485 0.3215 2.333 0.3745 ;
              RECT  1.9585 0.3215 2.0435 0.3745 ;
              RECT  1.6685 0.3215 1.7535 0.3745 ;
              RECT  1.3785 0.3215 1.4635 0.3745 ;
              RECT  1.0535 0.3215 1.138 0.3745 ;
              RECT  0.7635 0.3215 0.8485 0.3745 ;
              RECT  0.4735 0.3215 0.5585 0.3745 ;
              RECT  0.1835 0.3215 0.2685 0.364 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2825 0.53 0.728 0.5865 ;
              RECT  0.6715 0.502 0.728 0.5865 ;
              RECT  0.608 0.53 0.6645 0.6505 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3325 0.544 1.7995 0.601 ;
              RECT  1.4385 0.544 1.5305 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.012 0.544 3.0685 0.6505 ;
              RECT  2.9875 0.502 3.0295 0.5865 ;
              RECT  2.3475 0.544 3.0685 0.5865 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.362 0.445 3.811 0.502 ;
              RECT  3.362 0.445 3.5105 0.6325 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.384 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.384 0.042 ;
        END
    END VSS
END NOR4X8

MACRO AOI21X2
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.4415 1.1065 0.4985 ;
              RECT  1.032 0.3425 1.1065 0.4985 ;
              RECT  0.8765 0.4415 0.9615 0.523 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.417 0.6115 0.502 ;
              RECT  0.4665 0.417 0.523 0.516 ;
              RECT  0.1835 0.417 0.6115 0.4735 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.544 0.3955 0.636 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.852 0.5935 0.894 0.721 ;
              RECT  0.7635 0.5935 0.894 0.636 ;
              RECT  0.7635 0.2615 0.806 0.636 ;
              RECT  0.7495 0.304 0.806 0.516 ;
              RECT  0.4065 0.304 0.806 0.346 ;
              RECT  0.357 0.2895 0.4415 0.332 ;
        END
    END Y
END AOI21X2

MACRO DFFX4
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.881 0.403 3.2985 0.445 ;
              RECT  3.178 0.7175 3.2205 0.993 ;
              RECT  2.8705 0.7175 3.2205 0.76 ;
              RECT  2.8705 0.7175 2.9305 0.993 ;
              RECT  2.8705 0.5585 2.927 0.993 ;
              RECT  2.881 0.403 2.927 0.993 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.5985 0.7175 2.641 0.993 ;
              RECT  2.2165 0.311 2.6335 0.3535 ;
              RECT  2.3085 0.7175 2.641 0.76 ;
              RECT  2.319 0.311 2.3615 0.76 ;
              RECT  2.3085 0.424 2.351 0.993 ;
              RECT  2.305 0.424 2.3615 0.516 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.371 0.6645 0.7245 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.3995 0.1695 0.516 ;
              RECT  0.042 0.3995 0.0985 0.682 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END DFFX4

MACRO CLKBUFX12
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3575 0.6925 1.4 1.025 ;
              RECT  0.166 0.3355 1.4 0.378 ;
              RECT  1.3575 0.18 1.4 0.378 ;
              RECT  0.166 0.6925 1.4 0.735 ;
              RECT  1.0675 0.6925 1.11 1.025 ;
              RECT  1.0675 0.18 1.11 0.378 ;
              RECT  0.7775 0.6925 0.82 1.025 ;
              RECT  0.7775 0.18 0.82 0.378 ;
              RECT  0.4875 0.6925 0.53 1.025 ;
              RECT  0.4875 0.18 0.53 0.378 ;
              RECT  0.1835 0.6925 0.24 1.025 ;
              RECT  0.1975 0.18 0.24 0.378 ;
              RECT  0.166 0.3355 0.2085 0.735 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.562 1.7005 0.6185 ;
              RECT  1.598 0.562 1.6545 0.8695 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END CLKBUFX12

MACRO NOR2X2
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.357 0.629 0.806 0.6715 ;
              RECT  0.7495 0.5585 0.806 0.6715 ;
              RECT  0.7495 0.3885 0.7915 0.6715 ;
              RECT  0.212 0.3885 0.7915 0.431 ;
              RECT  0.502 0.332 0.544 0.431 ;
              RECT  0.357 0.629 0.3995 0.997 ;
              RECT  0.212 0.332 0.2545 0.431 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.629 0.286 0.6855 ;
              RECT  0.1835 0.629 0.24 0.9365 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.502 0.5935 0.5585 ;
              RECT  0.042 0.502 0.0985 0.6505 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END NOR2X2

MACRO TIELO
    CLASS CORE ;
    SIZE 0.424 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.113 0.0985 0.4665 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.424 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.424 0.042 ;
        END
    END VSS
END TIELO

MACRO SDFFHQX1
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0985 0.3815 0.141 1.0425 ;
              RECT  0.042 0.424 0.141 0.516 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.33 0.4415 3.3725 0.5265 ;
              RECT  2.782 0.456 3.3725 0.4985 ;
              RECT  3.277 0.4415 3.3725 0.4985 ;
              RECT  2.782 0.456 2.8245 0.668 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.0155 0.569 3.2595 0.6325 ;
              RECT  3.0155 0.569 3.2275 0.735 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.542 0.4595 2.5985 0.643 ;
              RECT  2.4465 0.4595 2.5985 0.516 ;
              RECT  2.4465 0.385 2.503 0.516 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3425 0.5515 0.3995 0.7315 ;
              RECT  0.325 0.5585 0.3815 0.887 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END SDFFHQX1

MACRO NOR3BX4
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.18 0.265 2.047 0.3075 ;
              RECT  1.5375 0.795 1.58 0.972 ;
              RECT  0.18 0.795 1.58 0.8375 ;
              RECT  0.654 0.795 0.6965 0.972 ;
              RECT  0.18 0.265 0.2225 0.8375 ;
              RECT  0.042 0.2895 0.2225 0.332 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.831 0.484 1.9195 0.5265 ;
              RECT  1.3715 0.569 1.8735 0.6115 ;
              RECT  1.831 0.484 1.8735 0.6115 ;
              RECT  1.3715 0.491 1.414 0.6115 ;
              RECT  1.064 0.491 1.414 0.5335 ;
              RECT  0.4665 0.569 1.1065 0.6115 ;
              RECT  1.064 0.491 1.1065 0.6115 ;
              RECT  0.4665 0.424 0.523 0.6115 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.135 0.502 2.22 0.5585 ;
              RECT  2.135 0.378 2.192 0.5585 ;
              RECT  1.9905 0.378 2.192 0.4985 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5305 0.456 1.6155 0.4985 ;
              RECT  1.5305 0.378 1.573 0.4985 ;
              RECT  0.951 0.378 1.573 0.4205 ;
              RECT  0.7315 0.456 0.993 0.4985 ;
              RECT  0.951 0.378 0.993 0.4985 ;
              RECT  0.7315 0.4415 0.8235 0.4985 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END NOR3BX4

MACRO INVX3
    CLASS CORE ;
    SIZE 0.5655 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.47 0.509 0.5265 0.5655 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.438 0.1235 0.5975 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.5655 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.5655 0.042 ;
        END
    END VSS
END INVX3

MACRO CLKXOR2X4
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.8165 0.5265 0.9015 ;
              RECT  0.484 0.2085 0.5265 0.293 ;
              RECT  0.4525 0.636 0.4945 0.859 ;
              RECT  0.1835 0.364 0.4945 0.4065 ;
              RECT  0.4525 0.251 0.4945 0.4065 ;
              RECT  0.1835 0.636 0.4945 0.6785 ;
              RECT  0.1835 0.5585 0.24 0.6785 ;
              RECT  0.1835 0.5585 0.2365 0.912 ;
              RECT  0.1835 0.3075 0.2365 0.4065 ;
              RECT  0.1835 0.3075 0.226 0.912 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.4345 1.6545 0.6505 ;
              RECT  1.3435 0.4345 1.6545 0.491 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6785 0.477 0.933 0.5335 ;
              RECT  0.6785 0.477 0.8235 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END CLKXOR2X4

MACRO DFFSRX1
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.728 0.742 0.7705 0.827 ;
              RECT  0.622 0.2825 0.7635 0.325 ;
              RECT  0.721 0.24 0.7635 0.325 ;
              RECT  0.608 0.742 0.7705 0.7845 ;
              RECT  0.608 0.6925 0.6645 0.7845 ;
              RECT  0.622 0.2825 0.6645 0.7845 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.912 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END QN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.5675 0.2895 4.624 0.3815 ;
              RECT  4.525 0.325 4.582 0.601 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1435 0.5585 4.2 0.654 ;
              RECT  4.016 0.5585 4.2 0.615 ;
              RECT  4.016 0.4275 4.0725 0.615 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7895 0.608 3.433 0.6505 ;
              RECT  2.7895 0.212 2.8315 0.6505 ;
              RECT  2.3365 0.212 2.8315 0.2545 ;
              RECT  1.6015 0.569 2.379 0.6115 ;
              RECT  2.3365 0.212 2.379 0.6115 ;
              RECT  2.287 0.4415 2.379 0.4985 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9085 0.509 1.0215 0.5655 ;
              RECT  0.735 0.576 0.965 0.6325 ;
              RECT  0.9085 0.509 0.965 0.6325 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END DFFSRX1

MACRO AO21X4
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.424 1.3715 0.516 ;
              RECT  1.1735 0.424 1.3715 0.4665 ;
              RECT  1.1735 0.318 1.216 0.753 ;
              RECT  1.156 0.714 1.1985 0.9895 ;
              RECT  0.866 0.601 1.216 0.643 ;
              RECT  0.721 0.318 1.216 0.3605 ;
              RECT  1.011 0.2615 1.0535 0.3605 ;
              RECT  0.866 0.601 0.9085 0.9895 ;
              RECT  0.721 0.2615 0.7635 0.3605 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.417 0.24 0.7705 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.3955 0.7705 ;
              RECT  0.339 0.431 0.3955 0.7705 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5585 0.537 0.7705 ;
              RECT  0.4805 0.431 0.537 0.7705 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END AO21X4

MACRO SDFFTRX2
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8625 0.5585 0.9475 0.6505 ;
              RECT  0.8625 0.403 0.9475 0.445 ;
              RECT  0.8625 0.403 0.905 0.912 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.403 0.523 0.516 ;
              RECT  0.4665 0.403 0.509 0.912 ;
              RECT  0.438 0.403 0.523 0.445 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.43 0.1905 4.4865 0.516 ;
              RECT  4.426 0.1555 4.483 0.247 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.267 0.7105 4.359 0.774 ;
              RECT  4.3025 0.456 4.359 0.774 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.963 0.5585 4.1965 0.615 ;
              RECT  3.963 0.5585 4.076 0.6325 ;
              RECT  3.963 0.456 4.0195 0.6325 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.012 0.5585 3.224 0.643 ;
              RECT  3.1675 0.484 3.224 0.643 ;
              RECT  3.012 0.5585 3.0685 0.682 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.424 1.23 0.7775 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END SDFFTRX2

MACRO SDFFX2
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4435 0.403 3.528 0.445 ;
              RECT  3.4645 0.403 3.507 0.958 ;
              RECT  3.4365 0.424 3.507 0.516 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.424 3.21 0.516 ;
              RECT  3.1535 0.403 3.196 0.958 ;
              RECT  3.111 0.403 3.196 0.445 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8705 0.325 2.927 0.6785 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.5585 0.9475 0.6505 ;
              RECT  0.834 0.5935 0.8905 0.8555 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.7035 0.523 0.919 ;
              RECT  0.311 0.7035 0.523 0.76 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.576 0.523 0.6325 ;
              RECT  0.1835 0.576 0.24 0.661 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END SDFFX2

MACRO NOR3X4
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.022 0.2895 2.0785 0.3815 ;
              RECT  0.647 0.795 2.0645 0.8375 ;
              RECT  2.022 0.265 2.0645 0.8375 ;
              RECT  0.18 0.265 2.0645 0.3075 ;
              RECT  1.5305 0.795 1.573 0.972 ;
              RECT  0.647 0.795 0.689 0.972 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.364 0.682 1.909 0.7245 ;
              RECT  1.8665 0.583 1.909 0.7245 ;
              RECT  1.078 0.6045 1.163 0.7245 ;
              RECT  0.0565 0.6715 0.4065 0.714 ;
              RECT  0.0565 0.5585 0.0985 0.714 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7465 0.424 1.796 0.5585 ;
              RECT  1.633 0.4735 1.796 0.516 ;
              RECT  1.739 0.424 1.796 0.516 ;
              RECT  1.2515 0.537 1.6755 0.5795 ;
              RECT  1.633 0.4735 1.6755 0.5795 ;
              RECT  1.2515 0.491 1.294 0.5795 ;
              RECT  0.965 0.491 1.294 0.5335 ;
              RECT  0.477 0.569 1.0075 0.6115 ;
              RECT  0.965 0.491 1.0075 0.6115 ;
              RECT  0.346 0.5585 0.5195 0.601 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4105 0.424 1.4955 0.4665 ;
              RECT  1.4105 0.378 1.453 0.4665 ;
              RECT  0.654 0.378 1.453 0.4205 ;
              RECT  0.59 0.4415 0.6965 0.4985 ;
              RECT  0.654 0.378 0.6965 0.4985 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END NOR3X4

MACRO AOI31X4
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3505 0.4345 2.5525 0.477 ;
              RECT  2.51 0.378 2.5525 0.477 ;
              RECT  2.4465 0.6925 2.503 0.7845 ;
              RECT  2.4465 0.4345 2.489 0.7845 ;
              RECT  2.411 0.7035 2.4535 0.788 ;
              RECT  2.082 0.7035 2.503 0.7455 ;
              RECT  2.22 0.378 2.2625 0.477 ;
              RECT  2.082 0.7035 2.1245 0.788 ;
              RECT  1.93 0.378 1.9725 0.477 ;
              RECT  1.64 0.378 1.6825 0.477 ;
              RECT  1.3505 0.378 1.393 0.477 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.576 0.5975 0.6325 ;
              RECT  0.3075 0.491 0.364 0.6325 ;
              RECT  0.272 0.491 0.364 0.548 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.852 0.569 1.177 0.6255 ;
              RECT  0.852 0.569 0.965 0.6325 ;
              RECT  0.852 0.491 0.9365 0.6325 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.0505 0.548 2.3755 0.6045 ;
              RECT  2.146 0.548 2.2375 0.6325 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.576 1.7925 0.6325 ;
        END
    END A2
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END AOI31X4

MACRO OAI32X2
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5025 0.3215 1.598 0.364 ;
              RECT  1.018 0.357 1.545 0.3995 ;
              RECT  1.3185 0.88 1.361 0.965 ;
              RECT  1.018 0.88 1.361 0.9225 ;
              RECT  1.223 0.3215 1.308 0.3995 ;
              RECT  1.018 0.357 1.0605 0.9225 ;
              RECT  0.5725 0.7245 1.0605 0.767 ;
              RECT  0.873 0.7105 1.0605 0.767 ;
              RECT  0.5725 0.7245 0.615 0.965 ;
        END
    END Y
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5975 0.537 0.654 ;
              RECT  0.325 0.5975 0.3815 0.795 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.47 0.82 0.555 ;
              RECT  0.608 0.47 0.6645 0.6505 ;
              RECT  0.332 0.47 0.82 0.5265 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.301 0.583 1.4845 0.6395 ;
              RECT  1.315 0.583 1.3715 0.8095 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.357 0.9475 0.516 ;
              RECT  0.166 0.357 0.9475 0.3995 ;
              RECT  0.166 0.357 0.2085 0.516 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.131 0.47 1.626 0.5125 ;
              RECT  1.1735 0.47 1.23 0.6505 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END OAI32X2

MACRO CLKXOR2X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0985 0.4735 0.141 0.912 ;
              RECT  0.042 0.424 0.1025 0.516 ;
              RECT  0.06 0.3675 0.1025 0.516 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.689 0.576 1.085 0.6185 ;
              RECT  0.873 0.576 0.965 0.6325 ;
              RECT  0.5655 0.59 0.7315 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.516 0.3815 0.8695 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END CLKXOR2X1

MACRO NOR4X6
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.164 0.636 3.2065 0.9685 ;
              RECT  2.874 0.6505 3.2065 0.6925 ;
              RECT  3.026 0.247 3.0685 0.516 ;
              RECT  3.012 0.41 3.0545 0.6925 ;
              RECT  0.233 0.41 3.0685 0.4525 ;
              RECT  2.874 0.6505 2.9165 0.8555 ;
              RECT  2.5385 0.7705 2.9165 0.813 ;
              RECT  2.7365 0.247 2.7785 0.4525 ;
              RECT  2.5385 0.6505 2.5805 0.8555 ;
              RECT  2.379 0.247 2.4215 0.4525 ;
              RECT  2.0895 0.247 2.1315 0.4525 ;
              RECT  1.7995 0.247 1.842 0.4525 ;
              RECT  1.4315 0.247 1.474 0.4525 ;
              RECT  1.1415 0.247 1.184 0.4525 ;
              RECT  0.813 0.247 0.8555 0.4525 ;
              RECT  0.523 0.247 0.5655 0.4525 ;
              RECT  0.233 0.247 0.2755 0.4525 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.523 0.523 0.6505 ;
              RECT  0.24 0.53 0.523 0.5865 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9825 0.537 1.2975 0.5935 ;
              RECT  1.0145 0.537 1.1135 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.523 2.22 0.6505 ;
              RECT  1.831 0.523 2.22 0.5795 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.616 0.523 2.9165 0.5795 ;
              RECT  2.7115 0.523 2.8035 0.6325 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END NOR4X6

MACRO AOI222X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.972 0.8485 1.23 0.8905 ;
              RECT  1.1735 0.6925 1.23 0.8905 ;
              RECT  1.1735 0.2895 1.216 0.8905 ;
              RECT  0.537 0.325 1.216 0.3675 ;
              RECT  1.025 0.2895 1.216 0.3675 ;
              RECT  0.972 0.8485 1.0145 0.933 ;
              RECT  0.537 0.2685 0.5795 0.3675 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4805 0.438 0.537 0.7775 ;
              RECT  0.4665 0.438 0.537 0.6505 ;
        END
    END B1
    PIN C1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.018 0.438 1.0885 0.7775 ;
        END
    END C1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.346 0.24 0.7 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.622 0.608 0.774 0.7775 ;
              RECT  0.608 0.5335 0.6645 0.6505 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8445 0.5585 0.9475 0.6505 ;
              RECT  0.8445 0.5585 0.9015 0.866 ;
        END
    END C0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.1555 0.385 0.5055 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END AOI222X1

MACRO NAND4X8
    CLASS CORE ;
    SIZE 4.2425 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.2275 0.403 4.1825 0.445 ;
              RECT  3.9735 0.668 4.016 0.9825 ;
              RECT  3.684 0.7035 4.016 0.7455 ;
              RECT  3.8605 0.403 3.917 0.516 ;
              RECT  3.8605 0.403 3.903 0.7455 ;
              RECT  3.684 0.7035 3.726 0.9825 ;
              RECT  2.234 0.721 3.726 0.7635 ;
              RECT  3.394 0.7035 3.4365 0.9825 ;
              RECT  3.104 0.668 3.1465 0.9825 ;
              RECT  2.814 0.721 2.8565 0.9825 ;
              RECT  2.524 0.668 2.5665 0.9825 ;
              RECT  2.234 0.668 2.2765 0.9825 ;
              RECT  1.6545 0.6855 2.2765 0.728 ;
              RECT  1.9445 0.668 1.9865 0.9825 ;
              RECT  1.6545 0.6855 1.697 0.9825 ;
              RECT  0.4945 0.721 1.697 0.7635 ;
              RECT  1.3645 0.721 1.407 0.9825 ;
              RECT  1.0745 0.668 1.117 0.9825 ;
              RECT  0.7845 0.721 0.827 0.9825 ;
              RECT  0.4945 0.6855 0.537 0.9825 ;
              RECT  0.205 0.7845 0.537 0.827 ;
              RECT  0.205 0.6855 0.247 0.9825 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.5585 0.728 0.6395 ;
              RECT  0.6715 0.555 0.728 0.6395 ;
              RECT  0.608 0.5585 0.6645 0.6505 ;
              RECT  0.2825 0.5585 0.728 0.615 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3185 0.5585 1.764 0.615 ;
              RECT  1.4565 0.5585 1.513 0.6505 ;
              RECT  1.3185 0.5585 1.513 0.6395 ;
              RECT  1.3185 0.555 1.375 0.6395 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.729 0.5585 2.786 0.6505 ;
              RECT  2.312 0.555 2.7715 0.5975 ;
              RECT  2.715 0.5125 2.7715 0.5975 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.3265 0.576 3.79 0.6325 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.2425 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.2425 0.042 ;
        END
    END VSS
END NAND4X8

MACRO SDFFSX4
    CLASS CORE ;
    SIZE 5.6565 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.416 0.5585 5.473 0.6505 ;
              RECT  5.3065 0.5585 5.473 0.601 ;
              RECT  5.3065 0.463 5.349 0.601 ;
              RECT  4.8895 0.463 5.349 0.5055 ;
              RECT  4.8895 0.463 4.932 0.728 ;
              RECT  4.8575 0.6855 4.9 0.7705 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.1155 0.576 5.236 0.7455 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.617 0.576 4.6735 0.813 ;
              RECT  4.5005 0.576 4.6735 0.6325 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.444 0.7035 4.5465 0.76 ;
              RECT  4.2 0.7105 4.5005 0.767 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.0935 0.2545 3.136 0.4735 ;
              RECT  2.8845 0.2545 3.136 0.2965 ;
              RECT  2.8845 0.2085 2.927 0.2965 ;
              RECT  2.1635 0.2085 2.927 0.251 ;
              RECT  2.1635 0.424 2.22 0.516 ;
              RECT  1.87 0.576 2.206 0.6185 ;
              RECT  2.1635 0.2085 2.206 0.6185 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.354 0.3815 1.3965 0.993 ;
              RECT  1.032 0.4735 1.3965 0.516 ;
              RECT  1.064 0.3815 1.1065 0.993 ;
              RECT  1.032 0.424 1.1065 0.516 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.3815 0.5265 0.912 ;
              RECT  0.1835 0.608 0.5265 0.6505 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
              RECT  0.1835 0.3815 0.2365 0.912 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.6565 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.6565 0.042 ;
        END
    END VSS
END SDFFSX4

MACRO DFFSHQX8
    CLASS CORE ;
    SIZE 4.384 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1505 0.636 4.3625 0.6925 ;
              RECT  4.267 0.4945 4.3625 0.6925 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.8675 0.576 4.08 0.6925 ;
              RECT  4.023 0.4945 4.08 0.6925 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.846 0.1905 2.8885 0.516 ;
              RECT  2.6905 0.1905 2.8885 0.233 ;
              RECT  2.022 0.166 2.7325 0.2085 ;
              RECT  2.022 0.2895 2.0785 0.3815 ;
              RECT  1.8275 0.562 2.0645 0.6045 ;
              RECT  2.022 0.166 2.0645 0.6045 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.926 0.3815 0.9685 0.951 ;
              RECT  0.042 0.424 0.9685 0.4665 ;
              RECT  0.636 0.3815 0.6785 0.951 ;
              RECT  0.346 0.3815 0.3885 0.951 ;
              RECT  0.0565 0.3815 0.0985 0.951 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.384 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.384 0.042 ;
        END
    END VSS
END DFFSHQX8

MACRO NOR4BX4
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7965 0.7035 2.839 0.8025 ;
              RECT  1.156 0.7035 2.839 0.7455 ;
              RECT  0.622 0.392 2.694 0.4345 ;
              RECT  2.6515 0.3355 2.694 0.4345 ;
              RECT  2.5065 0.7035 2.549 0.8025 ;
              RECT  2.3615 0.3355 2.404 0.4345 ;
              RECT  2.0715 0.3355 2.114 0.4345 ;
              RECT  1.7815 0.3355 1.824 0.4345 ;
              RECT  1.4915 0.3355 1.534 0.4345 ;
              RECT  1.156 0.7035 1.248 0.767 ;
              RECT  1.202 0.3355 1.2445 0.4345 ;
              RECT  1.156 0.392 1.1985 0.767 ;
              RECT  0.912 0.3355 0.9545 0.4345 ;
              RECT  0.622 0.3355 0.6645 0.4345 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1445 0.4595 0.2015 0.675 ;
              RECT  0.042 0.4595 0.2015 0.516 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.269 0.576 1.6225 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8345 0.576 2.227 0.6325 ;
              RECT  1.8345 0.5055 1.8915 0.6325 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4145 0.576 2.807 0.6325 ;
              RECT  2.4145 0.5055 2.471 0.6325 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END NOR4BX4

MACRO CLKINVX3
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.583 0.636 0.6255 0.912 ;
              RECT  0.293 0.438 0.6255 0.4805 ;
              RECT  0.583 0.3815 0.6255 0.4805 ;
              RECT  0.293 0.636 0.6255 0.6785 ;
              RECT  0.325 0.438 0.3815 0.6785 ;
              RECT  0.293 0.636 0.3355 0.912 ;
              RECT  0.293 0.3815 0.3355 0.4805 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5125 0.2225 0.668 ;
              RECT  0.166 0.438 0.2225 0.668 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END CLKINVX3

MACRO SDFFHQX4
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1815 0.463 3.652 0.5055 ;
              RECT  3.56 0.4415 3.652 0.5055 ;
              RECT  3.1815 0.463 3.224 0.615 ;
              RECT  3.1605 0.5725 3.203 0.6575 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.408 0.576 3.5775 0.6965 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.92 0.53 2.9765 0.6575 ;
              RECT  2.729 0.5935 2.9765 0.6505 ;
              RECT  2.729 0.5585 2.786 0.6505 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.4875 0.24 0.841 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.7175 0.753 0.76 ;
              RECT  0.7105 0.3815 0.753 0.76 ;
              RECT  0.371 0.3815 0.4135 0.601 ;
              RECT  0.325 0.5585 0.3815 0.76 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END SDFFHQX4

MACRO NOR3X6
    CLASS CORE ;
    SIZE 2.9695 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7315 0.8165 2.927 0.859 ;
              RECT  2.8845 0.385 2.927 0.859 ;
              RECT  2.8705 0.6925 2.927 0.859 ;
              RECT  2.6125 0.385 2.927 0.4275 ;
              RECT  2.6125 0.2085 2.655 0.4275 ;
              RECT  0.6185 0.251 2.655 0.293 ;
              RECT  2.4995 0.8165 2.542 0.9015 ;
              RECT  2.28 0.2085 2.3225 0.293 ;
              RECT  1.948 0.2085 1.9905 0.293 ;
              RECT  1.7285 0.8165 1.771 0.9015 ;
              RECT  1.6155 0.2085 1.658 0.4065 ;
              RECT  1.283 0.2085 1.3255 0.293 ;
              RECT  0.951 0.2085 0.993 0.293 ;
              RECT  0.7315 0.8165 0.774 0.9015 ;
              RECT  0.286 0.385 0.661 0.4275 ;
              RECT  0.6185 0.2085 0.661 0.4275 ;
              RECT  0.286 0.2085 0.3285 0.4275 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.761 0.537 2.8035 0.622 ;
              RECT  0.233 0.7035 2.8 0.7455 ;
              RECT  2.7575 0.5975 2.8 0.7455 ;
              RECT  2.008 0.6255 2.093 0.7455 ;
              RECT  1.1205 0.6255 1.2055 0.7455 ;
              RECT  0.233 0.576 0.2755 0.7455 ;
              RECT  0.166 0.576 0.2755 0.6325 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.59 2.683 0.6325 ;
              RECT  2.641 0.5125 2.683 0.6325 ;
              RECT  2.57 0.576 2.683 0.6325 ;
              RECT  2.1635 0.5125 2.206 0.6325 ;
              RECT  1.895 0.5125 2.206 0.555 ;
              RECT  1.276 0.59 1.937 0.6325 ;
              RECT  1.895 0.5125 1.937 0.6325 ;
              RECT  1.389 0.548 1.4315 0.6325 ;
              RECT  1.276 0.5125 1.3185 0.6325 ;
              RECT  1.0075 0.5125 1.3185 0.555 ;
              RECT  0.357 0.59 1.05 0.6325 ;
              RECT  1.0075 0.5125 1.05 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.2765 0.477 2.5205 0.5195 ;
              RECT  2.2765 0.3995 2.319 0.5195 ;
              RECT  1.7815 0.3995 2.319 0.4415 ;
              RECT  1.5025 0.477 1.824 0.5195 ;
              RECT  1.7815 0.3995 1.824 0.5195 ;
              RECT  1.5025 0.3995 1.545 0.5195 ;
              RECT  0.894 0.3995 1.545 0.4415 ;
              RECT  0.7315 0.456 0.9365 0.4985 ;
              RECT  0.894 0.3995 0.9365 0.4985 ;
              RECT  0.7315 0.4415 0.8235 0.4985 ;
              RECT  0.7315 0.4415 0.8165 0.5195 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.9695 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.9695 0.042 ;
        END
    END VSS
END NOR3X6

MACRO TLATNX1
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.188 0.279 2.245 0.912 ;
              RECT  2.146 0.3075 2.245 0.364 ;
              RECT  2.1705 0.279 2.245 0.364 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.3815 1.796 0.9475 ;
        END
    END QN
    PIN GN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.7105 1.5305 0.767 ;
              RECT  1.4385 0.5515 1.4955 0.8695 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.636 0.3745 0.6925 ;
              RECT  0.318 0.555 0.3745 0.6925 ;
              RECT  0.1835 0.555 0.24 0.6925 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END TLATNX1

MACRO AO21X2
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.894 0.424 0.9475 1.0465 ;
              RECT  0.8905 0.424 0.9475 0.516 ;
              RECT  0.8485 0.279 0.8905 0.4665 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.417 0.24 0.7705 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.378 0.325 0.4345 0.59 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.583 0.449 0.6645 0.7105 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END AO21X2

MACRO AOI31X2
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.064 0.668 1.1065 0.753 ;
              RECT  1.0465 0.194 1.0885 0.7105 ;
              RECT  1.032 0.424 1.0885 0.516 ;
              RECT  0.4945 0.2365 1.0885 0.279 ;
        END
    END Y
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5055 0.576 0.7455 0.661 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.265 0.463 0.7455 0.5055 ;
              RECT  0.325 0.463 0.3815 0.6505 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8165 0.424 0.9475 0.516 ;
              RECT  0.8165 0.35 0.859 0.516 ;
              RECT  0.152 0.35 0.859 0.392 ;
              RECT  0.152 0.35 0.194 0.491 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.35 1.3715 0.7035 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END AOI31X2

MACRO NOR3X2
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.226 1.0885 0.3815 ;
              RECT  0.601 0.721 1.0745 0.7635 ;
              RECT  1.032 0.226 1.0745 0.7635 ;
              RECT  0.173 0.226 1.0885 0.2685 ;
              RECT  0.601 0.721 0.643 0.806 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3425 0.5655 0.6505 0.622 ;
              RECT  0.3075 0.576 0.3995 0.6325 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.4525 0.8095 0.537 ;
              RECT  0.7495 0.4525 0.806 0.6505 ;
              RECT  0.339 0.4525 0.8095 0.4945 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.887 0.339 0.9295 0.4985 ;
              RECT  0.042 0.339 0.9295 0.3815 ;
              RECT  0.042 0.339 0.0985 0.516 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END NOR3X2

MACRO NOR3BX2
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.226 1.0605 0.2685 ;
              RECT  0.59 0.608 0.6325 0.933 ;
              RECT  0.042 0.608 0.6325 0.6505 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
              RECT  0.0565 0.226 0.0985 0.6505 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.5655 0.806 0.873 ;
              RECT  0.7035 0.5655 0.806 0.622 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.4525 0.9475 0.6505 ;
              RECT  0.403 0.4525 0.9475 0.4945 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.131 0.4525 1.23 0.6505 ;
              RECT  1.131 0.4525 1.1875 0.7635 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END NOR3BX2

MACRO DFFTRX1
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.2895 0.689 0.3745 ;
              RECT  0.636 0.629 0.6785 0.9475 ;
              RECT  0.622 0.2895 0.6645 0.6715 ;
              RECT  0.608 0.2895 0.6645 0.3815 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.912 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.258 3.21 0.6115 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.998 0.5195 3.0545 0.7105 ;
              RECT  2.8705 0.5585 3.0545 0.615 ;
              RECT  2.8705 0.5585 2.927 0.6505 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6925 0.9475 0.7495 ;
              RECT  0.8905 0.5515 0.9475 0.7495 ;
              RECT  0.7495 0.6925 0.806 0.7845 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END DFFTRX1

MACRO TLATXL
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.3355 2.22 0.7385 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5235 0.9615 1.6615 1.0535 ;
              RECT  1.605 0.286 1.6615 1.0535 ;
        END
    END QN
    PIN G
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.537 1.3715 0.8905 ;
        END
    END G
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.4525 0.7245 ;
              RECT  0.3955 0.4415 0.4525 0.7245 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END TLATXL

MACRO AO22X4
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.424 1.3715 0.516 ;
              RECT  1.315 0.346 1.3575 0.9225 ;
              RECT  1.025 0.647 1.3575 0.689 ;
              RECT  0.9295 0.346 1.3575 0.3885 ;
              RECT  1.191 0.332 1.276 0.3885 ;
              RECT  1.025 0.647 1.0675 0.9225 ;
              RECT  0.88 0.332 0.965 0.3745 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7315 0.7105 0.926 0.767 ;
              RECT  0.7315 0.576 0.7915 0.767 ;
              RECT  0.707 0.576 0.7915 0.6325 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3675 0.24 0.721 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.3675 0.523 0.721 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.3955 0.707 ;
              RECT  0.339 0.3675 0.3955 0.707 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END AO22X4

MACRO NAND4X6
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.012 0.424 3.3515 0.4665 ;
              RECT  3.309 0.247 3.3515 0.4665 ;
              RECT  3.164 0.636 3.2065 0.9685 ;
              RECT  2.874 0.721 3.2065 0.7635 ;
              RECT  3.012 0.5585 3.0685 0.6505 ;
              RECT  3.012 0.3675 3.0545 0.7635 ;
              RECT  2.7045 0.41 3.0545 0.4525 ;
              RECT  2.874 0.6505 2.9165 0.9685 ;
              RECT  2.5275 0.7705 2.9165 0.813 ;
              RECT  2.7045 0.3675 2.747 0.4525 ;
              RECT  2.5275 0.636 2.57 0.9685 ;
              RECT  2.2375 0.6715 2.57 0.714 ;
              RECT  2.2375 0.6715 2.28 0.9685 ;
              RECT  0.8835 0.721 2.28 0.7635 ;
              RECT  1.9055 0.6505 1.948 0.9685 ;
              RECT  1.6155 0.636 1.658 0.9685 ;
              RECT  1.2725 0.721 1.315 0.9685 ;
              RECT  0.8835 0.636 0.926 0.9685 ;
              RECT  0.304 0.7705 0.926 0.813 ;
              RECT  0.5935 0.636 0.636 0.9685 ;
              RECT  0.304 0.6505 0.346 0.9685 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.523 0.523 0.682 ;
              RECT  0.272 0.523 0.523 0.5795 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.544 1.4565 0.601 ;
              RECT  1.1735 0.523 1.23 0.6505 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.0045 0.544 2.188 0.601 ;
              RECT  2.1315 0.516 2.188 0.601 ;
              RECT  2.022 0.544 2.0785 0.6505 ;
              RECT  1.9335 0.523 2.061 0.5795 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.729 0.523 2.9415 0.5795 ;
              RECT  2.641 0.576 2.8035 0.6325 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END NAND4X6

MACRO SDFFSX2
    CLASS CORE ;
    SIZE 4.808 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.753 0.3815 0.8095 0.912 ;
              RECT  0.7495 0.424 0.8095 0.516 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.3815 0.24 0.912 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.3165 0.4415 4.5995 0.484 ;
              RECT  4.1645 0.456 4.5005 0.4985 ;
              RECT  4.3165 0.4135 4.359 0.4985 ;
              RECT  4.122 0.7245 4.207 0.767 ;
              RECT  4.1645 0.456 4.207 0.767 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4335 0.689 4.6735 0.7455 ;
              RECT  4.55 0.576 4.6735 0.7455 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.7225 0.3885 3.981 0.445 ;
              RECT  3.8605 0.3885 3.917 0.5405 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.56 0.7105 3.652 0.767 ;
              RECT  3.567 0.449 3.652 0.767 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3935 0.233 2.478 0.2755 ;
              RECT  2.1245 0.346 2.4355 0.3885 ;
              RECT  2.3935 0.233 2.4355 0.3885 ;
              RECT  2.1245 0.2225 2.167 0.3885 ;
              RECT  1.58 0.2225 2.167 0.265 ;
              RECT  1.3115 0.59 1.672 0.6325 ;
              RECT  1.58 0.576 1.672 0.6325 ;
              RECT  1.58 0.2225 1.6225 0.6325 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.808 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.808 0.042 ;
        END
    END VSS
END SDFFSX2

MACRO MX3X2
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.251 0.629 0.293 1.0465 ;
              RECT  0.251 0.2825 0.293 0.3675 ;
              RECT  0.219 0.325 0.2615 0.6715 ;
              RECT  0.166 0.4415 0.2615 0.4985 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7005 0.76 2.0785 0.8165 ;
              RECT  2.022 0.6925 2.0785 0.8165 ;
              RECT  1.7005 0.7245 1.757 0.8165 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8805 0.523 1.937 0.689 ;
              RECT  1.6935 0.523 1.937 0.5795 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3395 0.3675 1.3965 0.615 ;
              RECT  1.315 0.5585 1.3715 0.6965 ;
        END
    END B
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.3675 1.23 0.721 ;
        END
    END S1
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.364 0.7105 0.5585 0.767 ;
              RECT  0.502 0.5515 0.5585 0.767 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END MX3X2

MACRO NOR4X4
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.417 0.4205 2.489 0.463 ;
              RECT  2.4465 0.364 2.489 0.463 ;
              RECT  2.4075 0.7035 2.45 0.8025 ;
              RECT  0.7635 0.7035 2.45 0.7455 ;
              RECT  2.1565 0.364 2.199 0.463 ;
              RECT  2.1175 0.7035 2.16 0.8025 ;
              RECT  1.8665 0.364 1.909 0.463 ;
              RECT  1.5765 0.364 1.619 0.463 ;
              RECT  1.2865 0.364 1.329 0.463 ;
              RECT  0.997 0.364 1.039 0.463 ;
              RECT  0.7635 0.4205 0.806 0.7455 ;
              RECT  0.7495 0.5585 0.806 0.6505 ;
              RECT  0.707 0.364 0.7495 0.463 ;
              RECT  0.417 0.364 0.4595 0.463 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.247 0.615 0.6645 0.6715 ;
              RECT  0.608 0.5335 0.6645 0.6715 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.576 1.276 0.6325 ;
              RECT  1.2195 0.5335 1.276 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4915 0.576 1.817 0.6325 ;
              RECT  1.7215 0.548 1.817 0.6325 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.0045 0.576 2.418 0.6325 ;
              RECT  2.1955 0.548 2.252 0.6325 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END NOR4X4

MACRO OAI222XL
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.53 0.8695 1.202 0.912 ;
              RECT  1.1595 0.332 1.202 0.912 ;
              RECT  1.018 0.332 1.202 0.3745 ;
              RECT  1.032 0.8695 1.0995 1.0535 ;
              RECT  0.986 0.3215 1.0605 0.364 ;
              RECT  0.986 0.2155 1.0285 0.364 ;
              RECT  0.53 0.8695 0.5725 0.979 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.445 0.6645 0.799 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.445 0.24 0.799 ;
        END
    END A0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.431 0.9475 0.7845 ;
        END
    END C0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5405 0.385 0.6505 ;
              RECT  0.325 0.5405 0.3815 0.8905 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.445 1.0885 0.799 ;
        END
    END C1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.445 0.806 0.799 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OAI222XL

MACRO AOI222X4
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5955 0.7035 3.638 0.8025 ;
              RECT  1.347 0.7035 3.638 0.7455 ;
              RECT  3.3055 0.7035 3.348 0.8025 ;
              RECT  3.189 0.3355 3.3375 0.378 ;
              RECT  0.5865 0.35 3.224 0.392 ;
              RECT  3.0155 0.7035 3.058 0.8025 ;
              RECT  2.814 0.3355 2.899 0.392 ;
              RECT  2.7255 0.7035 2.768 0.8025 ;
              RECT  2.2695 0.3355 2.3545 0.392 ;
              RECT  1.658 0.3355 1.743 0.392 ;
              RECT  1.347 0.35 1.389 0.7455 ;
              RECT  1.2975 0.576 1.389 0.6325 ;
              RECT  0.9755 0.3355 1.0605 0.392 ;
              RECT  0.537 0.3355 0.622 0.378 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.743 0.576 2.2625 0.6325 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.449 0.576 1.0075 0.6325 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.867 0.576 3.3905 0.6325 ;
        END
    END C1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4915 0.463 2.5525 0.5055 ;
              RECT  1.58 0.576 1.672 0.6325 ;
              RECT  1.58 0.463 1.6225 0.6325 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.648 0.463 3.6415 0.5055 ;
              RECT  3.4185 0.4415 3.5105 0.5055 ;
        END
    END C0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2965 0.463 1.2265 0.5055 ;
              RECT  0.3075 0.4415 0.3995 0.5055 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END AOI222X4

MACRO CLKINVX6
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.781 0.636 0.8235 0.9685 ;
              RECT  0.2015 0.3285 0.8235 0.371 ;
              RECT  0.781 0.173 0.8235 0.371 ;
              RECT  0.491 0.636 0.8235 0.6785 ;
              RECT  0.608 0.5585 0.6645 0.6785 ;
              RECT  0.608 0.3285 0.6505 0.6785 ;
              RECT  0.491 0.636 0.5335 0.9685 ;
              RECT  0.491 0.173 0.5335 0.371 ;
              RECT  0.194 0.7705 0.5335 0.813 ;
              RECT  0.2015 0.173 0.2435 0.371 ;
              RECT  0.194 0.636 0.2365 0.9685 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1625 0.4415 0.516 0.4985 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END CLKINVX6

MACRO NOR4BBX2
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8805 0.424 1.937 0.516 ;
              RECT  1.8805 0.318 1.923 0.6115 ;
              RECT  1.863 0.569 1.9055 0.8095 ;
              RECT  1.2125 0.318 1.923 0.3605 ;
              RECT  1.7925 0.2615 1.8345 0.3605 ;
              RECT  1.5025 0.2615 1.545 0.3605 ;
              RECT  0.8905 0.2965 1.255 0.325 ;
              RECT  1.2125 0.2545 1.255 0.3605 ;
              RECT  0.94 0.318 1.923 0.339 ;
              RECT  0.8905 0.2825 0.9755 0.325 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.573 0.4595 1.81 0.516 ;
              RECT  1.573 0.4595 1.672 0.6325 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.5335 1.5025 0.654 ;
              RECT  1.446 0.431 1.5025 0.654 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2085 0.7105 0.4205 0.767 ;
              RECT  0.364 0.569 0.4205 0.767 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2085 0.4415 0.4205 0.4985 ;
              RECT  0.2085 0.4415 0.265 0.6395 ;
        END
    END BN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END NOR4BBX2

MACRO OR2X1
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.516 ;
              RECT  0.608 0.318 0.6505 0.6645 ;
              RECT  0.5935 0.2685 0.636 0.3535 ;
              RECT  0.59 0.6255 0.6325 0.912 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.304 0.576 0.424 0.6325 ;
              RECT  0.304 0.516 0.378 0.6325 ;
              RECT  0.304 0.516 0.3605 0.806 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0635 0.325 0.12 0.5865 ;
              RECT  0.042 0.2545 0.0985 0.3815 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END OR2X1

MACRO MX4X4
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5775 0.424 3.6345 0.516 ;
              RECT  2.959 0.424 3.6345 0.4665 ;
              RECT  3.4645 0.424 3.507 0.53 ;
              RECT  2.959 0.424 3.0015 0.509 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1145 0.576 3.394 0.6325 ;
              RECT  3.1145 0.576 3.171 0.707 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.45 0.7105 2.662 0.767 ;
              RECT  2.45 0.569 2.5065 0.767 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.287 0.569 2.379 0.788 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.3745 1.796 0.728 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.873 0.3075 0.9895 0.364 ;
              RECT  0.88 0.3075 0.9365 0.601 ;
        END
    END S1
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4845 0.6575 1.5695 0.7 ;
              RECT  1.4845 0.3285 1.5695 0.371 ;
              RECT  1.4845 0.3285 1.527 0.7 ;
              RECT  1.1735 0.608 1.527 0.6505 ;
              RECT  1.1525 0.6575 1.237 0.7 ;
              RECT  1.1735 0.608 1.237 0.7 ;
              RECT  1.1735 0.544 1.23 0.7 ;
              RECT  1.1735 0.3075 1.216 0.7 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END MX4X4

MACRO MDFFHQX1
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0985 0.3815 0.141 1.0425 ;
              RECT  0.042 0.424 0.141 0.516 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.33 0.4415 3.3725 0.5265 ;
              RECT  2.782 0.456 3.3725 0.4985 ;
              RECT  3.277 0.4415 3.3725 0.4985 ;
              RECT  2.782 0.456 2.8245 0.668 ;
        END
    END S0
    PIN D1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.0155 0.569 3.2595 0.6325 ;
              RECT  3.0155 0.569 3.2275 0.735 ;
        END
    END D1
    PIN D0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.542 0.4595 2.5985 0.643 ;
              RECT  2.4465 0.4595 2.5985 0.516 ;
              RECT  2.4465 0.385 2.503 0.516 ;
        END
    END D0
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3425 0.5515 0.3995 0.7315 ;
              RECT  0.325 0.5585 0.3815 0.887 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END MDFFHQX1

MACRO NOR4BX2
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.7035 1.7815 0.8025 ;
              RECT  0.9155 0.7035 1.7815 0.7455 ;
              RECT  0.6965 0.3425 1.6365 0.385 ;
              RECT  1.5945 0.286 1.6365 0.385 ;
              RECT  1.3045 0.286 1.347 0.385 ;
              RECT  0.986 0.286 1.0285 0.385 ;
              RECT  0.9155 0.3425 0.958 0.7455 ;
              RECT  0.8905 0.5585 0.958 0.6505 ;
              RECT  0.6965 0.286 0.7385 0.385 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.3215 0.615 ;
              RECT  0.2545 0.5195 0.3215 0.615 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0285 0.576 1.2515 0.6325 ;
              RECT  1.156 0.5655 1.2515 0.6325 ;
              RECT  1.0285 0.456 1.085 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.322 0.576 1.5555 0.6325 ;
              RECT  1.322 0.456 1.4385 0.6325 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.626 0.456 1.8135 0.6325 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END NOR4BX2

MACRO DFFSRHQX4
    CLASS CORE ;
    SIZE 5.2325 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.2135 0.905 3.68 0.9475 ;
              RECT  2.945 0.866 3.256 0.9085 ;
              RECT  2.379 0.951 2.9875 0.993 ;
              RECT  2.945 0.866 2.9875 0.993 ;
              RECT  2.379 0.7105 2.4215 0.993 ;
              RECT  2.1035 0.7105 2.4215 0.753 ;
              RECT  2.146 0.7105 2.2375 0.767 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.953 0.4415 5.211 0.5265 ;
              RECT  4.953 0.4415 5.0095 0.5935 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.437 0.576 4.656 0.668 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1345 0.4415 1.255 0.6115 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5975 0.293 0.6395 0.9475 ;
              RECT  0.3075 0.4735 0.6395 0.516 ;
              RECT  0.3075 0.424 0.3815 0.516 ;
              RECT  0.3075 0.293 0.35 0.9475 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.2325 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.2325 0.042 ;
        END
    END VSS
END DFFSRHQX4

MACRO NAND4BX2
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5695 0.3215 1.665 0.364 ;
              RECT  0.834 0.463 1.612 0.5055 ;
              RECT  1.5695 0.3215 1.612 0.5055 ;
              RECT  1.4955 0.788 1.559 0.986 ;
              RECT  0.6255 0.788 1.559 0.8305 ;
              RECT  1.2055 0.788 1.248 0.986 ;
              RECT  0.9155 0.788 0.958 0.986 ;
              RECT  0.8905 0.788 0.958 0.919 ;
              RECT  0.834 0.463 0.8765 0.8305 ;
              RECT  0.6255 0.788 0.668 0.986 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.127 0.576 0.2965 0.6325 ;
              RECT  0.127 0.4985 0.1835 0.6325 ;
              RECT  0.021 0.4985 0.1835 0.5585 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9475 0.576 1.1065 0.7175 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.177 0.601 1.446 0.7175 ;
              RECT  1.177 0.576 1.389 0.7175 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5165 0.629 1.817 0.6855 ;
              RECT  1.527 0.576 1.817 0.6855 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END NAND4BX2

MACRO AOI2BB1X4
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1235 0.3285 1.1985 0.371 ;
              RECT  1.156 0.272 1.1985 0.371 ;
              RECT  0.8695 0.8445 0.912 1.0425 ;
              RECT  0.866 0.272 0.9085 0.371 ;
              RECT  0.1235 0.8445 0.912 0.887 ;
              RECT  0.576 0.272 0.6185 0.371 ;
              RECT  0.431 0.8445 0.4735 1.0425 ;
              RECT  0.286 0.272 0.3285 0.371 ;
              RECT  0.166 0.8445 0.258 0.9015 ;
              RECT  0.1235 0.3285 0.166 0.887 ;
        END
    END Y
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.3075 1.3715 0.661 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.3535 1.6545 0.707 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2365 0.555 1.2405 0.5975 ;
              RECT  0.325 0.555 0.3815 0.6505 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END AOI2BB1X4

MACRO AO22X2
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0355 0.6925 1.0885 1.0465 ;
              RECT  1.032 0.293 1.0745 0.7845 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7245 0.675 0.806 0.7915 ;
              RECT  0.7245 0.463 0.781 0.7915 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.675 0.113 0.7845 ;
              RECT  0.0565 0.445 0.113 0.7845 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.4275 0.5405 0.7455 ;
              RECT  0.449 0.4275 0.5405 0.4985 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3215 0.576 0.378 0.7565 ;
              RECT  0.1835 0.576 0.378 0.6325 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END AO22X2

MACRO NOR4X2
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.714 0.9085 1.3715 0.951 ;
              RECT  1.329 0.3285 1.3715 0.951 ;
              RECT  1.315 0.827 1.3715 0.951 ;
              RECT  0.2435 0.3285 1.3715 0.371 ;
              RECT  1.1275 0.3145 1.2125 0.371 ;
              RECT  0.8165 0.3145 0.9015 0.371 ;
              RECT  0.5055 0.3145 0.59 0.371 ;
              RECT  0.194 0.3145 0.279 0.357 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.795 1.23 0.8375 ;
              RECT  1.1875 0.5795 1.23 0.8375 ;
              RECT  1.1735 0.6925 1.23 0.8375 ;
              RECT  0.1835 0.5795 0.226 0.8375 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.682 1.057 0.7245 ;
              RECT  1.0145 0.5975 1.057 0.7245 ;
              RECT  0.339 0.5585 0.3815 0.7245 ;
              RECT  0.325 0.5585 0.3815 0.6505 ;
              RECT  0.2965 0.59 0.3815 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9015 0.4415 1.1065 0.4985 ;
              RECT  0.4525 0.569 0.9435 0.6115 ;
              RECT  0.9015 0.4415 0.9435 0.6115 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4525 0.4415 0.806 0.4985 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END NOR4X2

MACRO DFFQX1
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.067 0.339 0.1235 1.018 ;
              RECT  0.042 0.424 0.1235 0.516 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.9515 0.7105 2.2415 0.767 ;
              RECT  1.9515 0.7105 2.0965 0.8305 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.509 0.3815 0.8625 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END DFFQX1

MACRO MX2XL
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.6925 1.0885 0.7845 ;
              RECT  1.032 0.1835 1.0745 0.979 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.5585 0.9475 0.6505 ;
              RECT  0.859 0.5935 0.9155 0.88 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.4065 0.7635 ;
              RECT  0.35 0.4345 0.4065 0.7635 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.477 0.7105 0.562 0.767 ;
              RECT  0.1975 0.834 0.5335 0.8905 ;
              RECT  0.477 0.7105 0.5335 0.8905 ;
              RECT  0.1975 0.6925 0.2545 0.8905 ;
              RECT  0.1835 0.6925 0.2545 0.7845 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END MX2XL

MACRO XOR2X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0985 0.4735 0.141 0.912 ;
              RECT  0.042 0.424 0.1025 0.516 ;
              RECT  0.06 0.3675 0.1025 0.516 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.689 0.576 1.085 0.6185 ;
              RECT  0.873 0.576 0.965 0.6325 ;
              RECT  0.5655 0.59 0.7315 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.516 0.3815 0.8695 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END XOR2X1

MACRO NAND4X4
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.941 0.371 2.6125 0.4135 ;
              RECT  2.57 0.3145 2.6125 0.4135 ;
              RECT  2.39 0.7035 2.432 0.965 ;
              RECT  0.7495 0.7035 2.432 0.7455 ;
              RECT  2.266 0.3145 2.3085 0.4135 ;
              RECT  2.1 0.7035 2.1425 0.965 ;
              RECT  0.7635 0.463 1.983 0.5055 ;
              RECT  1.941 0.371 1.983 0.5055 ;
              RECT  1.6935 0.7035 1.7355 0.965 ;
              RECT  1.4035 0.7035 1.446 0.965 ;
              RECT  1.0885 0.7035 1.131 0.965 ;
              RECT  0.799 0.7035 0.841 0.965 ;
              RECT  0.194 0.689 0.806 0.7315 ;
              RECT  0.7495 0.7035 0.841 0.7845 ;
              RECT  0.7635 0.463 0.806 0.7845 ;
              RECT  0.491 0.689 0.5335 0.965 ;
              RECT  0.194 0.689 0.2365 0.965 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1625 0.4415 0.516 0.4985 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.576 1.23 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.054 0.484 2.1385 0.5265 ;
              RECT  1.481 0.59 2.0965 0.6325 ;
              RECT  2.054 0.484 2.0965 0.6325 ;
              RECT  2.0045 0.576 2.0965 0.6325 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.45 0.484 2.5345 0.5405 ;
              RECT  2.1955 0.576 2.5065 0.6325 ;
              RECT  2.45 0.484 2.5065 0.6325 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END NAND4X4

MACRO AOI2BB1X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2615 0.293 0.346 0.3355 ;
              RECT  0.0565 0.3075 0.2965 0.35 ;
              RECT  0.1765 0.5335 0.219 1.0425 ;
              RECT  0.0565 0.5335 0.219 0.576 ;
              RECT  0.0565 0.3075 0.0985 0.576 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.5335 0.3955 0.7495 ;
              RECT  0.325 0.6925 0.3815 0.873 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5335 0.523 0.887 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6925 0.806 0.7845 ;
              RECT  0.707 0.4735 0.7635 0.7495 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END AOI2BB1X1

MACRO CLKINVX16
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.6575 2.1 0.7 ;
              RECT  2.0575 0.4135 2.1 0.7 ;
              RECT  2.022 0.6575 2.0785 0.7845 ;
              RECT  2.0255 0.6575 2.068 0.951 ;
              RECT  0.318 0.4135 2.1 0.456 ;
              RECT  2.0255 0.371 2.068 0.456 ;
              RECT  1.7145 0.403 1.7995 0.456 ;
              RECT  1.7355 0.6575 1.778 0.951 ;
              RECT  1.4245 0.403 1.5095 0.456 ;
              RECT  1.446 0.6575 1.488 0.951 ;
              RECT  1.1345 0.403 1.2195 0.456 ;
              RECT  1.156 0.6575 1.1985 0.951 ;
              RECT  0.286 0.7035 1.1985 0.7455 ;
              RECT  0.8445 0.403 0.9295 0.456 ;
              RECT  0.866 0.7035 0.9085 0.951 ;
              RECT  0.555 0.403 0.6395 0.456 ;
              RECT  0.576 0.7035 0.6325 0.951 ;
              RECT  0.265 0.403 0.35 0.445 ;
              RECT  0.286 0.7035 0.3285 0.951 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.364 0.544 1.9865 0.5865 ;
              RECT  0.449 0.544 0.5405 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END CLKINVX16

MACRO BUFX8
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.997 0.3885 1.092 0.431 ;
              RECT  1.0285 0.6575 1.071 0.972 ;
              RECT  0.159 0.3995 1.0285 0.4415 ;
              RECT  0.159 0.6575 1.071 0.7 ;
              RECT  0.7175 0.3885 0.8025 0.4415 ;
              RECT  0.7385 0.6575 0.781 0.972 ;
              RECT  0.4275 0.3885 0.5125 0.4415 ;
              RECT  0.449 0.6575 0.491 0.972 ;
              RECT  0.1835 0.3995 0.24 0.516 ;
              RECT  0.1835 0.3995 0.226 0.7 ;
              RECT  0.159 0.6575 0.2015 0.972 ;
              RECT  0.159 0.357 0.2015 0.4415 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4565 0.424 1.513 0.7775 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END BUFX8

MACRO AND2X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.615 0.3745 0.682 1.0465 ;
              RECT  0.5795 0.3745 0.682 0.4985 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.3885 0.8905 ;
              RECT  0.332 0.544 0.3885 0.8905 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0845 0.5655 0.141 0.8695 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END AND2X1

MACRO NAND4X2
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.226 0.9085 1.513 0.951 ;
              RECT  1.4565 0.827 1.513 0.951 ;
              RECT  1.4565 0.3285 1.499 0.951 ;
              RECT  0.8375 0.3285 1.499 0.371 ;
              RECT  1.223 0.9085 1.2655 0.993 ;
              RECT  0.8905 0.9085 0.933 0.993 ;
              RECT  0.7565 0.3145 0.873 0.357 ;
              RECT  0.5585 0.9085 0.601 0.993 ;
              RECT  0.226 0.9085 0.2685 0.993 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.795 1.3715 0.8375 ;
              RECT  1.315 0.5795 1.3715 0.8375 ;
              RECT  0.1835 0.5795 0.226 0.8375 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.682 1.1735 0.7245 ;
              RECT  1.131 0.5975 1.1735 0.7245 ;
              RECT  0.339 0.5585 0.3815 0.7245 ;
              RECT  0.325 0.5585 0.3815 0.6505 ;
              RECT  0.2965 0.59 0.3815 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.569 0.986 0.6115 ;
              RECT  0.9435 0.4415 0.986 0.6115 ;
              RECT  0.873 0.4415 0.986 0.4985 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.4415 0.8025 0.4985 ;
              RECT  0.608 0.2825 0.6645 0.4985 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END NAND4X2

MACRO DFFSRHQX1
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.3815 0.0985 0.912 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.267 0.576 4.359 0.6325 ;
              RECT  4.267 0.3145 4.3235 0.6325 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.652 0.576 3.9205 0.6325 ;
              RECT  3.652 0.576 3.7155 0.7105 ;
              RECT  3.652 0.569 3.7085 0.7105 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.602 0.9755 2.821 1.018 ;
              RECT  2.602 0.8625 2.6445 1.018 ;
              RECT  2.333 0.8625 2.6445 0.905 ;
              RECT  1.6225 0.9085 2.3755 0.951 ;
              RECT  2.333 0.8625 2.3755 0.951 ;
              RECT  1.6225 0.806 1.665 0.951 ;
              RECT  1.301 0.806 1.665 0.8485 ;
              RECT  1.032 0.8485 1.3435 0.8905 ;
              RECT  1.032 0.548 1.0885 0.6505 ;
              RECT  1.032 0.548 1.0745 0.8905 ;
              RECT  1.004 0.548 1.0885 0.59 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7315 0.576 0.933 0.6325 ;
              RECT  0.7315 0.502 0.788 0.6325 ;
              RECT  0.654 0.502 0.788 0.5585 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END DFFSRHQX1

MACRO TLATNTSCAX3
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4465 0.424 2.7785 0.4665 ;
              RECT  2.7365 0.3675 2.7785 0.4665 ;
              RECT  2.7045 0.636 2.747 0.912 ;
              RECT  2.4145 0.636 2.747 0.6785 ;
              RECT  2.4465 0.424 2.503 0.516 ;
              RECT  2.4465 0.3675 2.489 0.6785 ;
              RECT  2.4145 0.636 2.457 0.912 ;
        END
    END ECK
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.318 0.5405 0.654 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.318 0.3815 0.516 ;
              RECT  0.3075 0.424 0.364 0.654 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0245 0.371 0.1235 0.6325 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END TLATNTSCAX3

MACRO BUFX16
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.902 0.403 1.9975 0.445 ;
              RECT  1.9335 0.6395 1.976 0.951 ;
              RECT  0.1625 0.4135 1.9335 0.456 ;
              RECT  0.1625 0.6395 1.976 0.682 ;
              RECT  1.6225 0.403 1.7075 0.456 ;
              RECT  1.644 0.6395 1.686 0.951 ;
              RECT  1.3325 0.403 1.4175 0.456 ;
              RECT  1.354 0.6395 1.3965 0.951 ;
              RECT  1.0425 0.403 1.1275 0.456 ;
              RECT  1.064 0.6395 1.1065 0.951 ;
              RECT  0.753 0.403 0.8375 0.456 ;
              RECT  0.774 0.6395 0.8165 0.951 ;
              RECT  0.463 0.403 0.548 0.456 ;
              RECT  0.484 0.6395 0.5265 0.951 ;
              RECT  0.1835 0.6395 0.24 0.7845 ;
              RECT  0.1835 0.6395 0.2365 0.951 ;
              RECT  0.194 0.371 0.2365 0.456 ;
              RECT  0.1625 0.4135 0.205 0.682 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.576 2.6585 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END BUFX16

MACRO AOI33XL
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.025 0.827 1.0885 0.919 ;
              RECT  0.735 0.7845 1.0675 0.827 ;
              RECT  1.025 0.247 1.0675 0.919 ;
              RECT  0.569 0.247 1.0675 0.2895 ;
              RECT  0.735 0.7845 0.7775 0.894 ;
              RECT  0.569 0.205 0.6115 0.2895 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END A0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.424 0.523 0.7775 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.3605 0.82 0.445 ;
              RECT  0.7495 0.3605 0.806 0.7 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.3605 0.9475 0.714 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.1905 0.3955 0.4945 ;
              RECT  0.325 0.1555 0.3815 0.247 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.7775 ;
        END
    END B2
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END AOI33XL

MACRO TLATSRXL
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.654 0.346 0.7105 0.8625 ;
              RECT  0.608 0.424 0.7105 0.516 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.721 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4465 0.6925 2.595 0.7495 ;
              RECT  2.5385 0.576 2.595 0.7495 ;
              RECT  2.4465 0.6925 2.503 0.8375 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7215 0.576 1.8595 0.682 ;
              RECT  1.5555 0.576 1.8595 0.6325 ;
        END
    END RN
    PIN G
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.431 1.3715 0.7845 ;
        END
    END G
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.894 0.6785 1.131 0.7495 ;
              RECT  1.0145 0.576 1.131 0.7495 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END TLATSRXL

MACRO MXI2X8
    CLASS CORE ;
    SIZE 2.5455 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.326 0.6925 2.3685 1.0075 ;
              RECT  1.778 0.318 2.3685 0.3605 ;
              RECT  2.326 0.2755 2.3685 0.3605 ;
              RECT  1.4565 0.6925 2.3685 0.735 ;
              RECT  2.0575 0.3075 2.1 0.735 ;
              RECT  2.036 0.6925 2.0785 1.0075 ;
              RECT  2.015 0.3075 2.1 0.3605 ;
              RECT  1.725 0.3075 1.81 0.35 ;
              RECT  1.7465 0.6925 1.7885 1.0075 ;
              RECT  1.4565 0.6925 1.513 0.7845 ;
              RECT  1.4565 0.286 1.499 1.0075 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.4985 0.9475 0.852 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.456 0.4665 0.6505 ;
              RECT  0.325 0.456 0.3815 0.7245 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.795 0.5935 0.852 ;
              RECT  0.537 0.6115 0.5935 0.852 ;
              RECT  0.1975 0.7 0.2545 0.852 ;
              RECT  0.1835 0.6925 0.24 0.7845 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.5455 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.5455 0.042 ;
        END
    END VSS
END MXI2X8

MACRO CLKMX2X2
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.424 1.23 0.516 ;
              RECT  1.0605 0.424 1.23 0.4665 ;
              RECT  1.0605 0.3005 1.103 0.781 ;
              RECT  1.0355 0.7385 1.078 1.0145 ;
              RECT  1.0355 0.258 1.078 0.3425 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8625 0.576 0.9895 0.6325 ;
              RECT  0.8625 0.576 0.919 0.859 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.311 0.675 0.438 0.7315 ;
              RECT  0.325 0.449 0.3815 0.7315 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.8025 0.5655 0.859 ;
              RECT  0.509 0.6575 0.5655 0.859 ;
              RECT  0.1835 0.6925 0.24 0.859 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END CLKMX2X2

MACRO MX2X6
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7355 0.654 1.778 0.986 ;
              RECT  1.718 0.166 1.7605 0.385 ;
              RECT  1.704 0.3425 1.7465 0.6965 ;
              RECT  1.17 0.424 1.7465 0.4665 ;
              RECT  1.446 0.424 1.488 0.986 ;
              RECT  1.428 0.166 1.4705 0.4665 ;
              RECT  1.17 0.424 1.23 0.622 ;
              RECT  1.17 0.251 1.2125 0.622 ;
              RECT  1.156 0.5865 1.1985 0.986 ;
              RECT  1.138 0.2085 1.1805 0.293 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.477 0.9475 0.8305 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.4665 0.7035 ;
              RECT  0.41 0.4345 0.4665 0.7035 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.774 0.5935 0.8305 ;
              RECT  0.537 0.647 0.5935 0.8305 ;
              RECT  0.1835 0.647 0.2545 0.7845 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END MX2X6

MACRO MXI2X6
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.015 0.5585 2.0575 1.0465 ;
              RECT  2.015 0.205 2.0575 0.4875 ;
              RECT  1.983 0.445 2.0255 0.601 ;
              RECT  1.598 0.5585 2.0575 0.601 ;
              RECT  1.725 0.205 1.7675 1.0465 ;
              RECT  1.435 0.608 1.6545 0.6505 ;
              RECT  1.598 0.5585 1.6545 0.6505 ;
              RECT  1.598 0.4945 1.64 0.6505 ;
              RECT  1.435 0.4945 1.64 0.537 ;
              RECT  1.435 0.608 1.4775 1.0465 ;
              RECT  1.435 0.205 1.4775 0.537 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.537 0.9475 0.8905 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.4735 0.6505 ;
              RECT  0.417 0.516 0.4735 0.6505 ;
              RECT  0.325 0.5585 0.3815 0.7775 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.212 0.8485 0.5865 0.8905 ;
              RECT  0.544 0.6785 0.5865 0.8905 ;
              RECT  0.212 0.742 0.2545 0.8905 ;
              RECT  0.1835 0.6925 0.24 0.7845 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END MXI2X6

MACRO XOR3X1
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.287 0.576 2.379 0.661 ;
              RECT  2.287 0.47 2.3295 0.661 ;
              RECT  2.068 0.47 2.3295 0.5125 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.304 0.576 0.4525 0.6325 ;
              RECT  0.304 0.371 0.3605 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0635 0.4345 0.12 0.767 ;
              RECT  0.042 0.5585 0.12 0.6505 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.998 0.7245 3.0865 0.767 ;
              RECT  3.044 0.403 3.0865 0.767 ;
              RECT  2.9945 0.4415 3.0865 0.4985 ;
              RECT  2.998 0.403 3.0865 0.4985 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
END XOR3X1

MACRO MDFFHQX4
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1605 0.463 3.652 0.5055 ;
              RECT  3.56 0.4415 3.652 0.5055 ;
              RECT  3.1605 0.463 3.203 0.6575 ;
        END
    END S0
    PIN D1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.408 0.576 3.5775 0.6965 ;
        END
    END D1
    PIN D0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.92 0.53 2.9765 0.6575 ;
              RECT  2.729 0.5935 2.9765 0.6505 ;
              RECT  2.729 0.5585 2.786 0.6505 ;
        END
    END D0
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.4875 0.24 0.841 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.7175 0.753 0.76 ;
              RECT  0.7105 0.3815 0.753 0.76 ;
              RECT  0.371 0.3815 0.4135 0.601 ;
              RECT  0.325 0.5585 0.3815 0.76 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END MDFFHQX4

MACRO OAI211X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4415 0.827 0.827 0.8695 ;
              RECT  0.7845 0.311 0.827 0.8695 ;
              RECT  0.7495 0.827 0.806 1.025 ;
              RECT  0.7565 0.2685 0.799 0.3535 ;
              RECT  0.4415 0.827 0.484 1.025 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.636 0.205 0.767 ;
              RECT  0.148 0.537 0.205 0.767 ;
              RECT  0.042 0.636 0.0985 0.7845 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.4525 0.3815 0.7565 ;
              RECT  0.2755 0.4525 0.3815 0.509 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4525 0.5585 0.5585 0.6325 ;
              RECT  0.502 0.4525 0.5585 0.6325 ;
              RECT  0.4665 0.5585 0.523 0.7565 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.629 0.537 0.714 0.5935 ;
              RECT  0.629 0.2895 0.6855 0.5935 ;
              RECT  0.608 0.2895 0.6855 0.3815 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OAI211X1

MACRO TBUFXL
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.6925 1.2335 0.7845 ;
              RECT  1.191 0.3995 1.2335 0.7845 ;
              RECT  1.184 0.3425 1.2265 0.4275 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4415 0.2155 1.0005 0.258 ;
              RECT  0.272 0.682 0.5975 0.7245 ;
              RECT  0.555 0.4415 0.5975 0.7245 ;
              RECT  0.4415 0.4415 0.5975 0.484 ;
              RECT  0.4415 0.2155 0.484 0.484 ;
              RECT  0.3075 0.682 0.3995 0.767 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.141 0.555 0.484 0.6115 ;
              RECT  0.141 0.5265 0.24 0.6115 ;
              RECT  0.1835 0.424 0.24 0.6115 ;
        END
    END OE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END TBUFXL

MACRO DFFRX1
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6505 0.3075 0.6925 0.392 ;
              RECT  0.622 0.35 0.6645 1.0285 ;
              RECT  0.608 0.424 0.6645 0.516 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.912 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.269 0.569 1.534 0.6785 ;
              RECT  1.269 0.5335 1.389 0.6785 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.735 0.661 0.972 0.7495 ;
              RECT  0.735 0.576 0.965 0.7495 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.136 0.4415 3.2915 0.576 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END DFFRX1

MACRO AND3X1
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.332 0.9475 1.011 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.502 0.6645 0.8555 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3675 0.5585 0.424 0.6925 ;
              RECT  0.1835 0.5585 0.424 0.615 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.6925 0.113 0.827 ;
              RECT  0.0565 0.4875 0.113 0.827 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END AND3X1

MACRO OAI222X2
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.424 2.3615 0.516 ;
              RECT  0.4415 0.8165 2.3475 0.859 ;
              RECT  2.305 0.35 2.3475 0.859 ;
              RECT  1.7075 0.35 2.3475 0.392 ;
              RECT  1.9975 0.293 2.04 0.392 ;
              RECT  1.7815 0.8165 1.824 0.9015 ;
              RECT  1.7075 0.293 1.75 0.392 ;
              RECT  1.191 0.8165 1.2335 0.9015 ;
              RECT  0.4415 0.8165 0.484 0.9015 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.194 0.7035 0.6645 0.7455 ;
              RECT  0.608 0.5585 0.6645 0.7455 ;
              RECT  0.194 0.5975 0.2365 0.7455 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.7035 1.513 0.7455 ;
              RECT  1.4705 0.5975 1.513 0.7455 ;
              RECT  1.032 0.5585 1.0885 0.7455 ;
              RECT  1.004 0.59 1.0885 0.6325 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.022 0.5585 2.107 0.601 ;
              RECT  2.022 0.5585 2.0785 0.6505 ;
              RECT  1.598 0.7035 2.0645 0.7455 ;
              RECT  2.022 0.5585 2.0645 0.7455 ;
              RECT  1.598 0.5975 1.64 0.7455 ;
        END
    END C0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.477 0.4595 0.6325 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.711 0.548 1.9515 0.6325 ;
              RECT  1.895 0.463 1.9515 0.6325 ;
        END
    END C1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2975 0.463 1.4 0.6325 ;
              RECT  1.1595 0.463 1.4 0.5195 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END OAI222X2

MACRO OAI33X4
    CLASS CORE ;
    SIZE 4.101 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5885 0.3355 3.684 0.378 ;
              RECT  2.1425 0.371 3.6305 0.4135 ;
              RECT  3.309 0.3355 3.394 0.4135 ;
              RECT  3.019 0.3355 3.104 0.4135 ;
              RECT  2.729 0.3355 2.814 0.4135 ;
              RECT  2.6055 0.7035 2.648 0.8375 ;
              RECT  1.4315 0.7035 2.648 0.7455 ;
              RECT  2.4395 0.3355 2.524 0.4135 ;
              RECT  2.3085 0.7035 2.351 0.8375 ;
              RECT  2.1425 0.3355 2.227 0.4135 ;
              RECT  1.488 0.463 2.1845 0.5055 ;
              RECT  2.1425 0.3355 2.1845 0.5055 ;
              RECT  2.0185 0.7035 2.061 0.951 ;
              RECT  1.7215 0.7035 1.764 0.8375 ;
              RECT  1.488 0.463 1.5305 0.7455 ;
              RECT  1.4385 0.576 1.5305 0.6325 ;
              RECT  1.4315 0.7035 1.474 0.8375 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.429 0.576 3.7755 0.6325 ;
              RECT  3.429 0.484 3.486 0.6325 ;
        END
    END B0
    PIN B2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.22 0.576 2.5735 0.6325 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.463 1.23 0.6505 ;
              RECT  0.8835 0.576 1.23 0.6325 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.6015 0.576 1.955 0.6325 ;
        END
    END A2
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.35 0.5935 0.6645 0.6505 ;
              RECT  0.608 0.463 0.6645 0.6505 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.835 0.576 3.15 0.6325 ;
              RECT  2.835 0.484 2.945 0.6325 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.101 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.101 0.042 ;
        END
    END VSS
END OAI33X4

MACRO MXI2X4
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2515 0.304 1.6685 0.346 ;
              RECT  1.527 0.59 1.5695 0.9545 ;
              RECT  1.237 0.59 1.5695 0.6325 ;
              RECT  1.269 0.576 1.389 0.6325 ;
              RECT  1.347 0.304 1.389 0.6325 ;
              RECT  1.237 0.59 1.2795 0.9545 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.025 0.5655 1.0885 0.799 ;
              RECT  1.025 0.4525 1.0815 0.799 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.445 0.4525 0.502 0.6855 ;
              RECT  0.325 0.4525 0.502 0.6505 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5725 0.6965 0.841 0.7385 ;
              RECT  0.799 0.4205 0.841 0.7385 ;
              RECT  0.1975 0.7565 0.615 0.799 ;
              RECT  0.5725 0.654 0.615 0.799 ;
              RECT  0.1835 0.682 0.24 0.7845 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END MXI2X4

MACRO CLKAND2X4
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.163 0.668 1.23 0.9435 ;
              RECT  1.1735 0.5585 1.23 0.9435 ;
              RECT  1.1735 0.357 1.216 0.9435 ;
              RECT  0.8025 0.357 1.216 0.3995 ;
              RECT  0.873 0.668 1.23 0.7105 ;
              RECT  1.092 0.3005 1.1345 0.3995 ;
              RECT  0.873 0.668 0.9155 0.9435 ;
              RECT  0.8025 0.3005 0.8445 0.3995 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.187 0.576 0.5405 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2015 0.449 0.6185 0.5055 ;
              RECT  0.3075 0.4415 0.3995 0.5055 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END CLKAND2X4

MACRO DFFSX1
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.346 0.6645 0.912 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.159 0.3815 0.2155 0.912 ;
              RECT  0.042 0.424 0.2155 0.516 ;
        END
    END QN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.295 0.325 3.3515 0.6785 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.339 3.21 0.6925 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2975 0.576 1.5485 0.7 ;
              RECT  1.262 0.576 1.5485 0.6325 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END DFFSX1

MACRO FILL2
    CLASS CORE ;
    SIZE 0.2825 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.2825 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.2825 0.042 ;
        END
    END VSS
END FILL2

MACRO DFFNSRXL
    CLASS CORE ;
    SIZE 4.384 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.636 0.6325 0.6785 0.951 ;
              RECT  0.629 0.378 0.6715 0.463 ;
              RECT  0.608 0.5585 0.6645 0.668 ;
              RECT  0.622 0.4345 0.6645 0.668 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.3815 0.2225 0.721 ;
              RECT  0.042 0.424 0.2225 0.516 ;
        END
    END QN
    PIN CKN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.306 0.403 4.3625 0.6325 ;
              RECT  4.1825 0.403 4.3625 0.4985 ;
        END
    END CKN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.7545 0.424 3.811 0.689 ;
              RECT  3.712 0.378 3.7685 0.516 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.701 1.0145 3.065 1.057 ;
              RECT  2.701 0.8625 2.7435 1.057 ;
              RECT  1.347 0.8625 2.7435 0.905 ;
              RECT  1.347 0.636 1.4315 0.6785 ;
              RECT  1.347 0.636 1.389 0.905 ;
              RECT  1.2975 0.7105 1.389 0.767 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.873 0.6925 0.9295 0.8625 ;
              RECT  0.7495 0.6925 0.9295 0.7845 ;
              RECT  0.7495 0.6325 0.806 0.7845 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.384 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.384 0.042 ;
        END
    END VSS
END DFFNSRXL

MACRO OAI211X4
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.976 0.371 2.464 0.4135 ;
              RECT  2.4215 0.3145 2.464 0.4135 ;
              RECT  2.2765 0.7245 2.319 0.951 ;
              RECT  1.407 0.7245 2.319 0.767 ;
              RECT  2.1315 0.3145 2.174 0.4135 ;
              RECT  1.9865 0.7245 2.029 0.951 ;
              RECT  1.3715 0.463 2.0185 0.5055 ;
              RECT  1.976 0.371 2.0185 0.5055 ;
              RECT  1.697 0.7245 1.739 0.951 ;
              RECT  0.4945 0.7105 1.5305 0.753 ;
              RECT  1.407 0.7105 1.4495 0.951 ;
              RECT  1.3715 0.463 1.414 0.753 ;
              RECT  0.9615 0.7105 1.004 0.951 ;
              RECT  0.4945 0.7105 0.537 0.951 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4275 0.576 0.972 0.6325 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2155 0.463 1.191 0.5055 ;
              RECT  0.1835 0.4665 0.24 0.6505 ;
              RECT  0.1555 0.4665 0.24 0.509 ;
        END
    END A0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.5585 2.372 0.622 ;
              RECT  2.3155 0.537 2.372 0.622 ;
              RECT  2.1635 0.5585 2.22 0.6505 ;
              RECT  2.0715 0.5585 2.372 0.615 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4845 0.576 1.838 0.6325 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END OAI211X4

MACRO TLATNCAX8
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1605 0.371 3.203 0.986 ;
              RECT  2.291 0.6715 3.203 0.714 ;
              RECT  2.6125 0.4135 3.203 0.456 ;
              RECT  2.8495 0.403 2.934 0.456 ;
              RECT  2.8705 0.6715 2.913 0.986 ;
              RECT  2.5595 0.403 2.6445 0.445 ;
              RECT  2.5805 0.6715 2.623 0.986 ;
              RECT  2.291 0.424 2.3615 0.714 ;
              RECT  2.291 0.3815 2.333 0.986 ;
        END
    END ECK
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.378 0.7565 0.548 0.813 ;
              RECT  0.41 0.7105 0.548 0.813 ;
              RECT  0.41 0.5725 0.4665 0.813 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.134 0.7105 0.3075 0.767 ;
              RECT  0.251 0.53 0.3075 0.767 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END TLATNCAX8

MACRO BUFX12
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3575 0.6925 1.4 1.025 ;
              RECT  0.166 0.3355 1.4 0.378 ;
              RECT  1.3575 0.18 1.4 0.378 ;
              RECT  0.166 0.6925 1.4 0.735 ;
              RECT  1.0675 0.6925 1.11 1.025 ;
              RECT  1.0675 0.18 1.11 0.378 ;
              RECT  0.7775 0.6925 0.82 1.025 ;
              RECT  0.7775 0.18 0.82 0.378 ;
              RECT  0.4875 0.6925 0.53 1.025 ;
              RECT  0.4875 0.18 0.53 0.378 ;
              RECT  0.1835 0.6925 0.24 1.025 ;
              RECT  0.1975 0.18 0.24 0.378 ;
              RECT  0.166 0.3355 0.2085 0.735 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.562 1.7005 0.6185 ;
              RECT  1.598 0.562 1.6545 0.8695 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END BUFX12

MACRO SEDFFX1
    CLASS CORE ;
    SIZE 4.9495 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.6585 0.4415 2.701 0.774 ;
              RECT  2.57 0.4415 2.701 0.4985 ;
              RECT  2.57 0.3815 2.6125 0.4985 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.643 1.4 0.7 ;
              RECT  1.315 0.346 1.3715 0.7 ;
              RECT  1.276 0.346 1.3715 0.431 ;
        END
    END QN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.709 0.5585 4.8645 0.6925 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.438 2.3615 0.7915 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.6925 1.7285 0.7495 ;
              RECT  1.672 0.5125 1.7285 0.7495 ;
              RECT  1.598 0.6925 1.6545 0.7915 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3815 0.576 0.622 0.661 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.2365 1.0745 0.643 ;
              RECT  0.6255 0.2365 1.0745 0.279 ;
              RECT  0.6925 0.463 0.735 0.5515 ;
              RECT  0.2685 0.463 0.735 0.5055 ;
              RECT  0.6255 0.2365 0.668 0.5055 ;
              RECT  0.166 0.576 0.311 0.6325 ;
              RECT  0.2685 0.463 0.311 0.6325 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.9495 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.9495 0.042 ;
        END
    END VSS
END SEDFFX1

MACRO OAI33X2
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.008 0.7105 2.8495 0.753 ;
              RECT  2.807 0.668 2.8495 0.753 ;
              RECT  2.1425 0.7105 2.2375 0.767 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.7035 1.58 0.767 ;
              RECT  0.53 0.7035 1.58 0.7455 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.895 0.5975 2.7365 0.6395 ;
              RECT  1.8805 0.6925 1.937 0.7845 ;
              RECT  1.895 0.5975 1.937 0.7845 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.576 1.368 0.6325 ;
              RECT  0.3425 0.576 1.368 0.6185 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.484 2.623 0.5265 ;
              RECT  1.739 0.484 1.796 0.6505 ;
        END
    END B2
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2295 0.456 1.0605 0.4985 ;
              RECT  0.3075 0.4415 0.3995 0.4985 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9945 0.272 3.037 0.357 ;
              RECT  2.694 0.4065 3.005 0.449 ;
              RECT  2.9625 0.3145 3.005 0.449 ;
              RECT  0.59 0.8555 2.9625 0.898 ;
              RECT  2.92 0.4065 2.9625 0.898 ;
              RECT  2.683 0.293 2.768 0.3355 ;
              RECT  1.7925 0.371 2.7365 0.4135 ;
              RECT  2.683 0.293 2.7365 0.4135 ;
              RECT  2.372 0.293 2.457 0.4135 ;
              RECT  2.061 0.293 2.146 0.4135 ;
              RECT  1.7925 0.293 1.8345 0.4135 ;
              RECT  1.7215 0.3075 1.8345 0.364 ;
              RECT  1.75 0.293 1.8345 0.364 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END OAI33X2

MACRO EDFFHQX2
    CLASS CORE ;
    SIZE 3.6765 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.153 0.7495 2.245 0.806 ;
              RECT  2.153 0.3885 2.2375 0.445 ;
              RECT  2.153 0.3885 2.2095 0.806 ;
              RECT  2.022 0.5585 2.2095 0.6505 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4365 0.424 3.493 0.516 ;
              RECT  2.906 0.424 3.493 0.4665 ;
              RECT  2.9945 0.1975 3.037 0.4665 ;
              RECT  2.6795 0.1975 3.037 0.24 ;
              RECT  2.906 0.424 2.9485 0.5655 ;
              RECT  2.6795 0.1975 2.722 0.6925 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1465 0.537 3.3655 0.5935 ;
              RECT  3.1535 0.537 3.21 0.728 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.7105 0.3005 0.799 ;
              RECT  0.1625 0.5265 0.219 0.767 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.6765 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.6765 0.042 ;
        END
    END VSS
END EDFFHQX2

MACRO AND4X1
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.039 0.7105 1.1065 1.039 ;
              RECT  1.064 0.3995 1.1065 1.039 ;
              RECT  1.0075 0.3995 1.1065 0.4415 ;
              RECT  1.0075 0.357 1.05 0.4415 ;
              RECT  1.0145 0.7105 1.1065 0.767 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.767 0.548 0.8235 0.8835 ;
              RECT  0.7495 0.548 0.8235 0.6505 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5125 0.523 0.866 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.5125 0.3955 0.7495 ;
              RECT  0.325 0.6925 0.3815 0.852 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5125 0.24 0.8375 ;
              RECT  0.1555 0.537 0.24 0.5935 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END AND4X1

MACRO CLKMX2X8
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3085 0.35 2.351 1.0145 ;
              RECT  1.4385 0.7 2.351 0.742 ;
              RECT  1.7605 0.392 2.351 0.4345 ;
              RECT  1.9975 0.3815 2.082 0.4345 ;
              RECT  2.0185 0.7 2.061 1.0145 ;
              RECT  1.7075 0.3815 1.7925 0.424 ;
              RECT  1.7285 0.7 1.771 1.0145 ;
              RECT  1.4565 0.6925 1.513 0.7845 ;
              RECT  1.4565 0.3745 1.499 0.7845 ;
              RECT  1.4385 0.7 1.481 1.0145 ;
              RECT  1.414 0.3745 1.499 0.417 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.601 1.23 0.841 ;
              RECT  1.0605 0.601 1.23 0.6575 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.449 0.5055 0.5655 0.767 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.636 0.6115 0.721 0.654 ;
              RECT  0.3355 0.8375 0.6785 0.88 ;
              RECT  0.636 0.6115 0.6785 0.88 ;
              RECT  0.3355 0.675 0.378 0.88 ;
              RECT  0.1835 0.675 0.378 0.7845 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END CLKMX2X8

MACRO XNOR2X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.2895 0.2085 0.332 ;
              RECT  0.166 0.247 0.2085 0.332 ;
              RECT  0.0985 0.2895 0.141 0.9435 ;
              RECT  0.042 0.2895 0.141 0.3815 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0535 0.5195 1.138 0.576 ;
              RECT  0.841 0.576 1.11 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3745 0.3815 0.431 0.615 ;
              RECT  0.325 0.5585 0.3815 0.6855 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END XNOR2X1

MACRO AOI22X4
    CLASS CORE ;
    SIZE 2.5455 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.2555 0.7035 2.298 0.788 ;
              RECT  1.3855 0.7035 2.298 0.7455 ;
              RECT  1.884 0.3145 2.0325 0.357 ;
              RECT  1.9655 0.7035 2.008 0.788 ;
              RECT  0.5405 0.3285 1.9195 0.371 ;
              RECT  1.6755 0.7035 1.718 0.788 ;
              RECT  1.5095 0.3145 1.5945 0.371 ;
              RECT  1.3855 0.59 1.428 0.788 ;
              RECT  1.23 0.576 1.389 0.6325 ;
              RECT  1.23 0.3285 1.2725 0.6325 ;
              RECT  0.9295 0.3145 1.0145 0.371 ;
              RECT  0.491 0.3145 0.576 0.357 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5625 0.576 2.082 0.6325 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4415 0.576 0.9615 0.6325 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.463 1.1595 0.5265 ;
              RECT  1.117 0.4415 1.1595 0.5265 ;
              RECT  1.032 0.463 1.0885 0.6505 ;
              RECT  0.152 0.463 1.1595 0.5055 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3435 0.456 2.372 0.4985 ;
              RECT  1.4385 0.4415 1.5305 0.4985 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.5455 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.5455 0.042 ;
        END
    END VSS
END AOI22X4

MACRO SMDFFHQX4
    CLASS CORE ;
    SIZE 4.808 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4755 0.456 4.518 0.5405 ;
              RECT  4.4085 0.4415 4.5005 0.4985 ;
              RECT  3.9595 0.456 4.518 0.4985 ;
              RECT  3.9595 0.456 4.002 0.7 ;
        END
    END S0
    PIN D1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.193 0.569 4.405 0.6255 ;
              RECT  4.193 0.569 4.359 0.767 ;
        END
    END D1
    PIN D0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.719 0.3215 3.7755 0.675 ;
        END
    END D0
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5775 0.3215 3.6345 0.675 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.729 0.5585 2.9025 0.6505 ;
              RECT  2.846 0.4135 2.9025 0.6505 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.2965 0.24 0.6505 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.7 0.799 0.742 ;
              RECT  0.6645 0.378 0.707 0.502 ;
              RECT  0.6325 0.4595 0.675 0.742 ;
              RECT  0.325 0.5585 0.417 0.742 ;
              RECT  0.3745 0.378 0.417 0.742 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.808 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.808 0.042 ;
        END
    END VSS
END SMDFFHQX4

MACRO BUFX3
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4415 0.742 0.484 1.018 ;
              RECT  0.4135 0.2435 0.456 0.3285 ;
              RECT  0.152 0.742 0.484 0.7845 ;
              RECT  0.1235 0.3955 0.424 0.438 ;
              RECT  0.3815 0.286 0.424 0.438 ;
              RECT  0.1835 0.6925 0.24 0.7845 ;
              RECT  0.1835 0.3955 0.226 0.7845 ;
              RECT  0.152 0.742 0.194 1.018 ;
              RECT  0.1235 0.339 0.166 0.438 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.509 0.6645 0.8625 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END BUFX3

MACRO TLATNCAX20
    CLASS CORE ;
    SIZE 5.6565 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.494 0.555 5.5365 0.9895 ;
              RECT  5.473 0.251 5.515 0.4665 ;
              RECT  3.1535 0.555 5.5365 0.5975 ;
              RECT  5.441 0.424 5.4835 0.5975 ;
              RECT  5.204 0.555 5.2465 0.993 ;
              RECT  5.183 0.251 5.2255 0.5975 ;
              RECT  4.914 0.555 4.9565 0.993 ;
              RECT  4.893 0.251 4.9355 0.4665 ;
              RECT  4.861 0.424 4.9035 0.5975 ;
              RECT  4.624 0.555 4.6665 0.993 ;
              RECT  4.603 0.251 4.6455 0.5975 ;
              RECT  4.3345 0.555 4.3765 0.993 ;
              RECT  4.313 0.251 4.3555 0.484 ;
              RECT  4.2815 0.4415 4.3235 0.5975 ;
              RECT  4.0445 0.555 4.087 0.993 ;
              RECT  4.023 0.251 4.0655 0.5975 ;
              RECT  3.7545 0.555 3.797 0.993 ;
              RECT  3.7335 0.251 3.7755 0.4665 ;
              RECT  3.7015 0.424 3.744 0.5975 ;
              RECT  3.4645 0.555 3.507 0.993 ;
              RECT  3.4435 0.251 3.486 0.5975 ;
              RECT  3.1745 0.555 3.217 0.993 ;
              RECT  3.1535 0.251 3.196 0.6505 ;
        END
    END ECK
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.24 0.7845 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.6565 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.6565 0.042 ;
        END
    END VSS
END TLATNCAX20

MACRO AOI22X2
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.011 0.781 1.3435 0.8235 ;
              RECT  1.301 0.7035 1.3435 0.8235 ;
              RECT  0.502 0.293 1.191 0.3355 ;
              RECT  1.011 0.59 1.0535 0.8235 ;
              RECT  0.7315 0.59 1.0535 0.6325 ;
              RECT  0.7315 0.576 0.866 0.6325 ;
              RECT  0.8235 0.293 0.866 0.6325 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.463 0.5055 0.5265 0.6785 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.523 1.23 0.728 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.301 0.576 1.5305 0.6325 ;
              RECT  1.301 0.41 1.3855 0.6325 ;
              RECT  1.0605 0.41 1.3855 0.4525 ;
              RECT  0.9365 0.463 1.103 0.5055 ;
              RECT  1.0605 0.41 1.103 0.5055 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5935 0.449 0.753 0.5055 ;
              RECT  0.339 0.4065 0.6505 0.463 ;
              RECT  0.166 0.4415 0.3955 0.4985 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END AOI22X2

MACRO MXI3X4
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.428 0.332 1.8455 0.3745 ;
              RECT  1.7145 0.332 1.757 0.9545 ;
              RECT  1.4565 0.608 1.757 0.6505 ;
              RECT  1.4565 0.5585 1.513 0.6505 ;
              RECT  1.4565 0.5585 1.499 0.7245 ;
              RECT  1.4245 0.682 1.467 0.9545 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.121 0.456 2.623 0.4985 ;
              RECT  2.287 0.4415 2.379 0.4985 ;
              RECT  2.287 0.4415 2.351 0.5405 ;
              RECT  2.121 0.456 2.1635 0.7175 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3545 0.6115 2.6655 0.668 ;
              RECT  2.57 0.569 2.6655 0.668 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8805 0.445 1.937 0.799 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9545 0.6325 1.039 0.675 ;
              RECT  0.9545 0.502 0.997 0.675 ;
              RECT  0.728 0.502 0.997 0.544 ;
              RECT  0.728 0.484 0.806 0.544 ;
              RECT  0.7495 0.424 0.806 0.544 ;
              RECT  0.5405 0.544 0.7705 0.5865 ;
              RECT  0.4985 0.5585 0.583 0.601 ;
        END
    END S1
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1235 0.325 0.18 0.562 ;
              RECT  0.042 0.325 0.18 0.3815 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END MXI3X4

MACRO TLATNCAX2
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4735 0.4805 0.53 0.721 ;
              RECT  0.4665 0.3675 0.523 0.516 ;
        END
    END ECK
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.849 0.576 1.9865 0.661 ;
              RECT  1.849 0.4735 1.9055 0.7455 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.424 0.3815 0.516 ;
              RECT  0.2685 0.4595 0.325 0.721 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END TLATNCAX2

MACRO OAI2BB1X2
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5655 0.7845 0.608 1.0465 ;
              RECT  0.042 0.7845 0.608 0.827 ;
              RECT  0.12 0.431 0.463 0.4735 ;
              RECT  0.4205 0.3745 0.463 0.4735 ;
              RECT  0.2755 0.7845 0.318 1.0465 ;
              RECT  0.042 0.6925 0.1625 0.827 ;
              RECT  0.12 0.431 0.1625 0.827 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.233 0.544 0.6505 0.601 ;
              RECT  0.325 0.544 0.3815 0.6505 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.767 0.544 0.972 0.601 ;
              RECT  0.767 0.4415 0.8235 0.601 ;
              RECT  0.721 0.4415 0.8235 0.4985 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.827 1.23 0.919 ;
              RECT  1.156 0.583 1.2125 0.8835 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OAI2BB1X2

MACRO MXI2X2
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.424 1.3715 0.516 ;
              RECT  1.315 0.3815 1.3575 0.9435 ;
              RECT  1.3045 0.325 1.347 0.424 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.4945 1.149 0.6505 ;
              RECT  1.032 0.4945 1.0885 0.788 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.311 0.5585 0.5405 0.675 ;
              RECT  0.484 0.4945 0.5405 0.675 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6115 0.5935 0.8485 0.636 ;
              RECT  0.806 0.4945 0.8485 0.636 ;
              RECT  0.1975 0.7455 0.654 0.788 ;
              RECT  0.6115 0.5935 0.654 0.788 ;
              RECT  0.1835 0.6715 0.24 0.7845 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END MXI2X2

MACRO FILL64
    CLASS CORE ;
    SIZE 9.0505 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 9.0505 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 9.0505 0.042 ;
        END
    END VSS
END FILL64

MACRO SMDFFHQX1
    CLASS CORE ;
    SIZE 4.2425 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.06 0.3815 0.1025 0.9475 ;
              RECT  0.042 0.424 0.1025 0.516 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.0515 0.456 4.094 0.5405 ;
              RECT  3.5885 0.456 4.094 0.4985 ;
              RECT  3.7015 0.4415 3.7935 0.4985 ;
              RECT  3.5355 0.544 3.6305 0.5865 ;
              RECT  3.5885 0.456 3.6305 0.5865 ;
              RECT  3.5355 0.544 3.5775 0.735 ;
        END
    END S0
    PIN D1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.924 0.569 3.981 0.767 ;
              RECT  3.7685 0.569 3.981 0.654 ;
        END
    END D1
    PIN D0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.295 0.3425 3.3515 0.6965 ;
        END
    END D0
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.424 3.21 0.7775 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4995 0.424 2.556 0.714 ;
              RECT  2.4465 0.4135 2.503 0.5795 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.6505 0.3605 0.707 ;
              RECT  0.304 0.5515 0.3605 0.707 ;
              RECT  0.1835 0.6505 0.24 0.7845 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.2425 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.2425 0.042 ;
        END
    END VSS
END SMDFFHQX1

MACRO TLATSRX2
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.0545 0.5585 3.21 0.6505 ;
              RECT  3.0545 0.3955 3.097 0.661 ;
              RECT  3.0225 0.6185 3.065 0.951 ;
              RECT  3.0225 0.3535 3.065 0.438 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.57 0.4415 2.662 0.4985 ;
              RECT  2.457 0.4415 2.662 0.484 ;
              RECT  2.457 0.3355 2.4995 0.643 ;
              RECT  2.443 0.601 2.485 0.951 ;
              RECT  2.443 0.293 2.485 0.378 ;
        END
    END QN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.146 0.7105 2.3225 0.767 ;
              RECT  2.146 0.562 2.2305 0.767 ;
              RECT  2.146 0.562 2.2025 0.795 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.6395 1.3715 0.7845 ;
              RECT  1.1065 0.6395 1.3715 0.6965 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.438 0.4665 0.4945 0.707 ;
              RECT  0.325 0.4665 0.4945 0.6505 ;
        END
    END D
    PIN G
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.3745 1.6545 0.728 ;
        END
    END G
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END TLATSRX2

MACRO INVX20
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4995 0.509 2.556 0.5655 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.509 0.106 0.615 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END INVX20

MACRO AOI32X4
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.899 0.7035 2.9415 0.788 ;
              RECT  2.029 0.7035 2.9415 0.7455 ;
              RECT  0.59 0.2365 2.7185 0.279 ;
              RECT  2.609 0.7035 2.6515 0.788 ;
              RECT  2.319 0.7035 2.3615 0.788 ;
              RECT  2.029 0.576 2.0965 0.788 ;
              RECT  1.8665 0.576 2.0965 0.6325 ;
              RECT  1.8665 0.2365 1.909 0.6325 ;
        END
    END Y
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7845 0.654 1.354 0.6965 ;
              RECT  1.3115 0.576 1.354 0.6965 ;
              RECT  0.7845 0.59 0.827 0.6965 ;
              RECT  0.6045 0.576 0.8235 0.6325 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.206 0.576 2.7255 0.6325 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.184 0.463 1.64 0.5055 ;
              RECT  0.898 0.5405 1.2265 0.583 ;
              RECT  1.184 0.463 1.2265 0.583 ;
              RECT  0.898 0.463 0.94 0.583 ;
              RECT  0.378 0.463 0.94 0.5055 ;
              RECT  0.4665 0.463 0.523 0.6505 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.424 1.796 0.516 ;
              RECT  1.739 0.35 1.7815 0.516 ;
              RECT  1.711 0.463 1.796 0.5055 ;
              RECT  0.265 0.35 1.7815 0.392 ;
              RECT  1.011 0.35 1.096 0.47 ;
              RECT  0.265 0.35 0.3075 0.491 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.9795 0.456 3.0155 0.4985 ;
              RECT  1.9795 0.4415 2.2375 0.4985 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END AOI32X4

MACRO SDFFQX1
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.3815 0.0985 0.9475 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.485 0.456 2.945 0.4985 ;
              RECT  2.6055 0.4415 2.945 0.4985 ;
              RECT  2.6055 0.4135 2.648 0.4985 ;
              RECT  2.485 0.456 2.5275 0.569 ;
              RECT  2.4675 0.5265 2.51 0.7105 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7115 0.569 2.9765 0.6255 ;
              RECT  2.7115 0.569 2.8035 0.714 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.227 0.438 2.2835 0.7105 ;
              RECT  2.146 0.4415 2.2835 0.4985 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.6505 0.357 0.707 ;
              RECT  0.3005 0.5515 0.357 0.707 ;
              RECT  0.1835 0.6505 0.24 0.788 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END SDFFQX1

MACRO INVX4
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.615 0.445 0.6715 0.5655 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.509 0.106 0.615 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END INVX4

MACRO CLKMX2X12
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3155 0.6505 2.358 1.0465 ;
              RECT  2.2835 0.212 2.326 0.6925 ;
              RECT  1.156 0.5585 2.326 0.601 ;
              RECT  2.0255 0.5585 2.068 1.0465 ;
              RECT  1.994 0.212 2.036 0.601 ;
              RECT  1.7355 0.5585 1.778 1.0465 ;
              RECT  1.704 0.212 1.7465 0.601 ;
              RECT  1.446 0.5585 1.488 1.0465 ;
              RECT  1.414 0.212 1.4565 0.601 ;
              RECT  1.156 0.5585 1.23 0.6505 ;
              RECT  1.156 0.3355 1.1985 1.0465 ;
              RECT  1.0885 0.3355 1.1985 0.378 ;
              RECT  1.0885 0.293 1.131 0.378 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.562 0.9475 0.7845 ;
              RECT  0.866 0.7 0.9225 0.8905 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.4805 0.3955 0.7635 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.7315 0.569 0.788 ;
              RECT  0.1835 0.834 0.523 0.8905 ;
              RECT  0.4665 0.7315 0.523 0.8905 ;
              RECT  0.1835 0.6505 0.24 0.8905 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END CLKMX2X12

MACRO DFFSRXL
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6645 0.364 0.707 0.449 ;
              RECT  0.6255 0.4065 0.668 0.9295 ;
              RECT  0.608 0.424 0.668 0.516 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.3815 0.2225 0.721 ;
              RECT  0.042 0.424 0.2225 0.516 ;
        END
    END QN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.426 0.5335 4.483 0.887 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.002 0.5585 4.101 0.654 ;
              RECT  4.002 0.3425 4.0585 0.654 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.648 0.5655 3.256 0.608 ;
              RECT  2.648 0.212 2.6905 0.608 ;
              RECT  2.1955 0.212 2.6905 0.2545 ;
              RECT  1.442 0.4985 2.2375 0.5405 ;
              RECT  2.1955 0.212 2.2375 0.5405 ;
              RECT  2.146 0.4415 2.2375 0.5405 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7385 0.7105 0.965 0.82 ;
              RECT  0.8445 0.636 0.965 0.82 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END DFFSRXL

MACRO EDFFHQX8
    CLASS CORE ;
    SIZE 4.808 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1425 0.424 3.1815 0.4665 ;
              RECT  3.1395 0.3815 3.1815 0.4665 ;
              RECT  2.1175 0.682 3.072 0.7245 ;
              RECT  2.807 0.3815 2.8495 0.4665 ;
              RECT  2.4745 0.3815 2.517 0.4665 ;
              RECT  2.1635 0.5585 2.22 0.7245 ;
              RECT  2.1775 0.424 2.22 0.7245 ;
              RECT  2.1425 0.3815 2.1845 0.4665 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4155 0.4415 4.642 0.5055 ;
              RECT  4.1825 0.456 4.642 0.4985 ;
              RECT  4.2705 0.2295 4.313 0.4985 ;
              RECT  3.956 0.2295 4.313 0.272 ;
              RECT  3.956 0.2295 3.9985 0.6325 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.2955 0.576 4.649 0.6325 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.537 0.24 0.8905 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.808 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.808 0.042 ;
        END
    END VSS
END EDFFHQX8

MACRO MXI3X2
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4495 0.403 1.534 0.4595 ;
              RECT  1.4565 0.403 1.513 0.9435 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4285 0.4415 2.5205 0.4985 ;
              RECT  2.4285 0.346 2.5135 0.4985 ;
              RECT  1.902 0.346 2.5135 0.3885 ;
              RECT  2.0505 0.346 2.093 0.4805 ;
              RECT  1.902 0.346 1.9445 0.636 ;
              RECT  1.863 0.5935 1.9055 0.6785 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.5585 2.358 0.675 ;
              RECT  2.3015 0.4595 2.358 0.675 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.6225 0.3215 1.679 0.615 ;
              RECT  1.598 0.5585 1.6545 0.6505 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.509 0.7105 1.092 0.753 ;
              RECT  1.05 0.615 1.092 0.753 ;
              RECT  0.8625 0.502 0.905 0.753 ;
              RECT  0.59 0.7105 0.682 0.767 ;
              RECT  0.509 0.622 0.5515 0.753 ;
        END
    END S1
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.6925 0.1835 0.7495 ;
              RECT  0.127 0.516 0.1835 0.7495 ;
              RECT  0.042 0.6925 0.0985 0.7845 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END MXI3X2

MACRO MX2X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0465 0.6925 1.23 0.7845 ;
              RECT  1.0465 0.2615 1.0885 1.0005 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.873 0.509 0.965 0.7705 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.449 0.7175 ;
              RECT  0.392 0.431 0.449 0.7175 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.788 0.576 0.8445 ;
              RECT  0.5195 0.59 0.576 0.8445 ;
              RECT  0.1835 0.6925 0.24 0.8445 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END MX2X1

MACRO SEDFFHQX4
    CLASS CORE ;
    SIZE 5.798 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.593 0.4415 5.6355 0.5265 ;
              RECT  4.999 0.456 5.6355 0.4985 ;
              RECT  5.3985 0.4415 5.6355 0.4985 ;
              RECT  4.9565 0.5865 5.0415 0.629 ;
              RECT  4.999 0.456 5.0415 0.629 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.2255 0.569 5.5225 0.6255 ;
              RECT  5.2255 0.569 5.349 0.682 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.536 0.576 4.7725 0.6645 ;
              RECT  4.536 0.491 4.5925 0.6645 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.719 0.502 3.7755 0.8555 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.592 0.502 3.6485 0.682 ;
              RECT  3.4185 0.548 3.6485 0.6325 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.3815 0.5265 0.9545 ;
              RECT  0.1835 0.4735 0.5265 0.516 ;
              RECT  0.1835 0.424 0.24 0.516 ;
              RECT  0.1835 0.3815 0.2365 0.9545 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.798 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.798 0.042 ;
        END
    END VSS
END SEDFFHQX4

MACRO MXI4X4
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4185 0.576 3.68 0.6185 ;
              RECT  3.27 0.774 3.5105 0.8165 ;
              RECT  3.468 0.576 3.5105 0.8165 ;
              RECT  3.4185 0.576 3.5105 0.6325 ;
              RECT  2.0045 0.887 3.3125 0.9295 ;
              RECT  3.27 0.774 3.3125 0.9295 ;
              RECT  2.0045 0.548 2.047 0.9295 ;
        END
    END S1
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8845 0.4135 3.422 0.456 ;
              RECT  3.3795 0.265 3.422 0.456 ;
              RECT  3.1675 0.661 3.302 0.7035 ;
              RECT  3.1675 0.4135 3.21 0.7035 ;
              RECT  3.1535 0.4135 3.21 0.516 ;
              RECT  2.8845 0.661 2.9695 0.7035 ;
              RECT  2.927 0.4135 2.9695 0.7035 ;
              RECT  2.8845 0.265 2.927 0.456 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.6925 1.8205 0.8485 ;
              RECT  1.7285 0.53 1.785 0.7775 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.6925 1.2445 0.8485 ;
              RECT  1.1875 0.509 1.2445 0.8485 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0465 0.509 1.103 0.7775 ;
              RECT  1.032 0.6925 1.0885 0.8485 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6115 0.41 0.852 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5725 0.484 0.629 0.6645 ;
              RECT  0.1835 0.484 0.629 0.5405 ;
              RECT  0.1835 0.484 0.24 0.6505 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END MXI4X4

MACRO DLY1X4
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3045 0.636 1.347 0.912 ;
              RECT  1.0145 0.424 1.347 0.4665 ;
              RECT  1.3045 0.3675 1.347 0.4665 ;
              RECT  1.0145 0.636 1.347 0.6785 ;
              RECT  1.032 0.5585 1.0885 0.6785 ;
              RECT  1.032 0.424 1.0745 0.6785 ;
              RECT  1.0145 0.636 1.057 0.912 ;
              RECT  1.0145 0.3675 1.057 0.4665 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.548 0.3145 0.6325 ;
              RECT  0.166 0.548 0.2225 0.8095 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END DLY1X4

MACRO SDFFSRHQX2
    CLASS CORE ;
    SIZE 5.798 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3145 0.827 0.3815 0.919 ;
              RECT  0.3145 0.728 0.357 0.919 ;
              RECT  0.2825 0.523 0.325 0.7705 ;
              RECT  0.2545 0.3815 0.2965 0.5655 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.5575 0.5055 5.614 0.6505 ;
              RECT  4.9495 0.463 5.6 0.5055 ;
              RECT  4.9495 0.463 4.992 0.661 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.257 0.576 5.487 0.7175 ;
              RECT  5.218 0.601 5.487 0.6575 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.709 0.3535 4.7655 0.707 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.3945 0.576 4.6385 0.6325 ;
              RECT  4.582 0.4665 4.6385 0.6325 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7435 0.905 3.2805 0.9475 ;
              RECT  2.7435 0.8165 2.786 0.9475 ;
              RECT  2.4745 0.8165 2.786 0.859 ;
              RECT  1.909 0.912 2.517 0.9545 ;
              RECT  2.4745 0.8165 2.517 0.9545 ;
              RECT  1.909 0.6645 1.9515 0.9545 ;
              RECT  1.216 0.6645 1.9515 0.707 ;
              RECT  1.216 0.576 1.2585 0.707 ;
              RECT  1.156 0.576 1.2585 0.6325 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.852 0.53 1.085 0.5865 ;
              RECT  0.8905 0.53 0.9475 0.707 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.798 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.798 0.042 ;
        END
    END VSS
END SDFFSRHQX2

MACRO XOR2XL
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0845 0.311 0.141 0.834 ;
              RECT  0.042 0.424 0.141 0.516 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6185 0.576 1.0885 0.6185 ;
              RECT  0.799 0.5655 0.8835 0.6185 ;
              RECT  0.7315 0.576 0.8235 0.6325 ;
              RECT  0.6185 0.576 0.661 0.661 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.378 0.583 0.4345 0.7495 ;
              RECT  0.325 0.6925 0.3815 0.8835 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END XOR2XL

MACRO SEDFFHQX1
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.4735 2.549 0.516 ;
              RECT  2.5065 0.3815 2.549 0.516 ;
              RECT  2.464 0.4735 2.5065 0.912 ;
              RECT  2.305 0.424 2.3615 0.516 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.426 0.431 4.483 0.7845 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.0045 0.576 2.1035 0.7 ;
              RECT  1.9125 0.576 2.1035 0.6325 ;
              RECT  1.9125 0.4805 1.9975 0.6325 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2195 0.4415 1.276 0.6645 ;
              RECT  1.0885 0.4415 1.276 0.4985 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3355 0.5585 0.523 0.6855 ;
              RECT  0.3355 0.463 0.392 0.6855 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.636 0.35 0.6785 0.491 ;
              RECT  0.2225 0.35 0.6785 0.392 ;
              RECT  0.2225 0.35 0.265 0.484 ;
              RECT  0.166 0.4415 0.258 0.4985 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END SEDFFHQX1

MACRO TLATNXL
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.286 2.22 0.721 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.894 1.665 0.979 ;
              RECT  1.598 0.286 1.6545 0.979 ;
        END
    END QN
    PIN GN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4565 0.537 1.513 0.8905 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.675 0.339 0.7845 ;
              RECT  0.2825 0.537 0.339 0.7845 ;
              RECT  0.1835 0.675 0.24 0.7915 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END TLATNXL

MACRO OAI2BB2XL
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.813 1.3435 0.8555 ;
              RECT  1.301 0.251 1.3435 0.8555 ;
              RECT  1.0995 0.859 1.248 0.9015 ;
              RECT  1.156 0.813 1.248 0.9015 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4565 0.424 1.513 0.516 ;
              RECT  1.414 0.4595 1.4705 0.735 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.3885 1.23 0.742 ;
        END
    END B1
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.417 0.3815 0.7705 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3535 0.24 0.707 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END OAI2BB2XL

MACRO OR4XL
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.2615 1.0885 0.9295 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.477 0.4595 0.5335 0.767 ;
              RECT  0.4665 0.424 0.523 0.516 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.3955 0.7845 ;
              RECT  0.339 0.445 0.3955 0.7845 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END D
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7915 0.417 0.8485 0.728 ;
              RECT  0.7495 0.417 0.8485 0.516 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END OR4XL

MACRO FILL8
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END FILL8

MACRO DFFQXL
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.35 0.0985 0.926 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.948 0.5975 2.1 0.654 ;
              RECT  1.93 0.781 2.0965 0.8375 ;
              RECT  1.948 0.5975 2.0965 0.8375 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1695 0.6925 0.3425 0.8375 ;
              RECT  0.286 0.601 0.3425 0.8375 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END DFFQXL

MACRO AND2XL
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.615 0.3745 0.6645 0.873 ;
              RECT  0.608 0.424 0.6645 0.516 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.827 0.523 0.997 ;
              RECT  0.4415 0.668 0.4985 0.8835 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.258 0.615 ;
              RECT  0.2015 0.53 0.258 0.615 ;
              RECT  0.042 0.5585 0.0985 0.7245 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END AND2XL

MACRO CLKBUFX3
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4415 0.742 0.484 1.018 ;
              RECT  0.4135 0.2435 0.456 0.3285 ;
              RECT  0.152 0.742 0.484 0.7845 ;
              RECT  0.1235 0.3955 0.424 0.438 ;
              RECT  0.3815 0.286 0.424 0.438 ;
              RECT  0.1835 0.6925 0.24 0.7845 ;
              RECT  0.1835 0.3955 0.226 0.7845 ;
              RECT  0.152 0.742 0.194 1.018 ;
              RECT  0.1235 0.339 0.166 0.438 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.509 0.6645 0.8625 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END CLKBUFX3

MACRO DFFTRXL
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6325 0.371 0.689 0.456 ;
              RECT  0.622 0.636 0.6785 0.827 ;
              RECT  0.608 0.403 0.6645 0.6925 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.721 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.033 0.325 3.09 0.622 ;
              RECT  3.012 0.2895 3.0685 0.3815 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8705 0.53 2.9625 0.5865 ;
              RECT  2.8705 0.2685 2.927 0.5865 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6575 0.919 0.714 ;
              RECT  0.8625 0.629 0.919 0.714 ;
              RECT  0.7495 0.6575 0.806 0.919 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END DFFTRXL

MACRO OR2X2
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.516 ;
              RECT  0.5405 0.6395 0.6505 0.682 ;
              RECT  0.608 0.3145 0.6505 0.682 ;
              RECT  0.5405 0.3145 0.6505 0.357 ;
              RECT  0.5405 0.6395 0.583 0.972 ;
              RECT  0.5405 0.272 0.583 0.357 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2895 0.576 0.424 0.6325 ;
              RECT  0.2895 0.576 0.364 0.8165 ;
              RECT  0.2895 0.5405 0.346 0.8165 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.325 0.106 0.636 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OR2X2

MACRO DLY2X4
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.5935 1.513 0.76 ;
              RECT  1.4565 0.424 1.513 0.76 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.548 0.788 0.59 0.9435 ;
              RECT  0.548 0.251 0.59 0.3355 ;
              RECT  0.516 0.293 0.5585 0.8305 ;
              RECT  0.258 0.424 0.5585 0.4665 ;
              RECT  0.258 0.424 0.3815 0.516 ;
              RECT  0.258 0.35 0.3005 0.9435 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END DLY2X4

MACRO NAND2X1
    CLASS CORE ;
    SIZE 0.424 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3355 0.537 0.392 0.636 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.067 0.569 0.152 0.6925 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2085 0.4345 0.265 0.5265 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.424 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.424 0.042 ;
        END
    END VSS
END NAND2X1

MACRO MXI4X2
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.2845 0.5585 3.3515 0.6505 ;
              RECT  3.2845 0.3995 3.341 0.7245 ;
              RECT  3.256 0.3995 3.341 0.456 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1205 0.7105 1.3575 0.8835 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4595 0.4595 0.516 0.608 ;
              RECT  0.1835 0.4595 0.516 0.516 ;
              RECT  0.1835 0.4595 0.2435 0.6505 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.813 0.7175 1.05 0.8835 ;
              RECT  0.813 0.7105 0.965 0.8835 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6785 0.516 0.735 ;
              RECT  0.325 0.5865 0.3815 0.806 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.507 0.59 3.652 0.6325 ;
              RECT  3.56 0.5405 3.652 0.6325 ;
              RECT  2.3365 0.887 3.5495 0.9295 ;
              RECT  3.507 0.59 3.5495 0.9295 ;
              RECT  2.3365 0.6185 2.4395 0.661 ;
              RECT  2.397 0.5585 2.4395 0.661 ;
              RECT  2.3365 0.6185 2.379 0.9295 ;
        END
    END S1
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.022 0.438 2.0785 0.7915 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END MXI4X2

MACRO AOI32X2
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.513 0.781 1.5555 0.866 ;
              RECT  1.223 0.781 1.5555 0.8235 ;
              RECT  0.576 0.3075 1.4315 0.35 ;
              RECT  1.223 0.7105 1.2655 0.866 ;
              RECT  1.0145 0.7105 1.2655 0.753 ;
              RECT  1.0145 0.7105 1.1065 0.767 ;
              RECT  1.064 0.3075 1.1065 0.767 ;
        END
    END Y
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3675 0.647 0.6045 0.7035 ;
              RECT  0.3075 0.7105 0.424 0.767 ;
              RECT  0.3675 0.647 0.424 0.767 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.5335 0.806 0.6505 ;
              RECT  0.3675 0.5335 0.806 0.576 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.336 0.6185 1.6545 0.7105 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.4205 0.9475 0.5795 ;
              RECT  0.2545 0.4205 0.9475 0.463 ;
              RECT  0.2545 0.4205 0.2965 0.5795 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7075 0.4415 1.7925 0.5655 ;
              RECT  1.177 0.4415 1.7925 0.4985 ;
              RECT  1.177 0.4415 1.2655 0.5655 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END AOI32X2

MACRO DFFNSRX2
    CLASS CORE ;
    SIZE 4.9495 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.5675 0.6925 4.624 0.7845 ;
              RECT  4.4935 0.6925 4.624 0.7495 ;
              RECT  4.4935 0.3815 4.55 0.7495 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1435 0.3815 4.2 0.7845 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.3955 0.8905 ;
              RECT  0.325 0.5515 0.3815 0.8905 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.516 2.22 0.6785 ;
              RECT  2.082 0.516 2.22 0.6505 ;
              RECT  2.082 0.4065 2.1385 0.6505 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8275 0.576 2.0115 0.6325 ;
              RECT  1.8275 0.4065 1.884 0.6325 ;
        END
    END SN
    PIN CKN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.5585 0.2545 0.8905 ;
              RECT  0.1835 0.5515 0.24 0.6505 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.9495 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.9495 0.042 ;
        END
    END VSS
END DFFNSRX2

MACRO OR3X4
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.424 1.23 0.516 ;
              RECT  1.011 0.424 1.23 0.4665 ;
              RECT  0.9295 0.7565 1.0535 0.799 ;
              RECT  1.011 0.2965 1.0535 0.799 ;
              RECT  0.9685 0.2545 1.011 0.339 ;
              RECT  0.6395 0.643 1.0535 0.6855 ;
              RECT  0.9295 0.7565 0.972 1.032 ;
              RECT  0.6965 0.2965 1.0535 0.339 ;
              RECT  0.647 0.2825 0.7315 0.325 ;
              RECT  0.6395 0.643 0.682 1.032 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.523 0.523 0.8765 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.226 0.4735 0.2825 0.7495 ;
              RECT  0.1835 0.6925 0.24 0.7845 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.431 0.0985 0.7845 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OR3X4

MACRO DFFRXL
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.583 0.35 0.707 0.392 ;
              RECT  0.6645 0.3075 0.707 0.392 ;
              RECT  0.583 0.6925 0.6645 0.7845 ;
              RECT  0.583 0.35 0.6255 0.8625 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.148 0.3815 0.205 0.721 ;
              RECT  0.042 0.424 0.205 0.516 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.262 0.509 1.5025 0.6785 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.873 0.576 0.965 0.6325 ;
              RECT  0.873 0.576 0.9295 0.894 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.136 0.4415 3.2915 0.576 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END DFFRXL

MACRO FILL16
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END FILL16

MACRO XOR3XL
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.287 0.576 2.379 0.661 ;
              RECT  2.287 0.47 2.3295 0.661 ;
              RECT  2.068 0.47 2.3295 0.5125 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.7105 0.403 0.767 ;
              RECT  0.3075 0.4525 0.364 0.767 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.067 0.4595 0.1235 0.788 ;
              RECT  0.042 0.5585 0.1235 0.6505 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.998 0.735 3.0865 0.7775 ;
              RECT  3.044 0.403 3.0865 0.7775 ;
              RECT  2.9945 0.4415 3.0865 0.4985 ;
              RECT  2.998 0.403 3.0865 0.4985 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
END XOR3XL

MACRO CLKBUFX6
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.403 1.0885 0.7565 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.629 0.647 0.6715 0.9685 ;
              RECT  0.042 0.4205 0.6715 0.463 ;
              RECT  0.629 0.247 0.6715 0.463 ;
              RECT  0.042 0.647 0.6715 0.689 ;
              RECT  0.339 0.647 0.3815 0.9685 ;
              RECT  0.339 0.247 0.3815 0.463 ;
              RECT  0.042 0.5585 0.0985 0.689 ;
              RECT  0.042 0.247 0.0915 0.9685 ;
        END
    END Y
END CLKBUFX6

MACRO AOI222XL
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.2895 1.3715 0.3815 ;
              RECT  1.1205 0.714 1.3575 0.7565 ;
              RECT  1.315 0.1905 1.3575 0.7565 ;
              RECT  0.5935 0.1905 1.3575 0.233 ;
              RECT  1.1205 0.714 1.163 0.8445 ;
              RECT  0.5935 0.1695 0.636 0.2545 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.59 0.576 0.774 0.6325 ;
              RECT  0.59 0.4065 0.7245 0.6325 ;
        END
    END B1
    PIN C1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1455 0.5865 1.2445 0.643 ;
              RECT  1.1735 0.332 1.23 0.643 ;
        END
    END C1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0245 0.576 0.2365 0.6325 ;
              RECT  0.152 0.4345 0.2365 0.6325 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.424 0.9475 0.7315 ;
              RECT  0.8445 0.5265 0.9475 0.583 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.018 0.304 1.0885 0.516 ;
              RECT  1.018 0.304 1.0745 0.643 ;
        END
    END C0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.576 0.41 0.6325 ;
              RECT  0.3075 0.325 0.392 0.6325 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END AOI222XL

MACRO OR4X6
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4775 0.371 2.1 0.4135 ;
              RECT  2.0575 0.194 2.1 0.4135 ;
              RECT  1.994 0.742 2.036 0.9685 ;
              RECT  1.704 0.742 2.036 0.7845 ;
              RECT  1.704 0.6925 1.937 0.7845 ;
              RECT  1.8805 0.371 1.923 0.7845 ;
              RECT  1.7675 0.194 1.81 0.4135 ;
              RECT  1.704 0.6925 1.7465 0.9685 ;
              RECT  1.414 0.6925 1.937 0.735 ;
              RECT  1.4775 0.194 1.52 0.4135 ;
              RECT  1.414 0.6925 1.4565 0.9685 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.6925 1.23 0.7845 ;
              RECT  0.212 0.827 1.216 0.8695 ;
              RECT  1.1735 0.569 1.216 0.8695 ;
              RECT  0.212 0.629 0.2545 0.8695 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.714 1.103 0.7565 ;
              RECT  1.0605 0.629 1.103 0.7565 ;
              RECT  0.325 0.6505 0.41 0.7565 ;
              RECT  0.325 0.5585 0.3815 0.7565 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4805 0.601 0.965 0.643 ;
              RECT  0.9225 0.4415 0.965 0.643 ;
              RECT  0.873 0.4415 0.965 0.4985 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4805 0.4735 0.8025 0.53 ;
              RECT  0.4805 0.4415 0.682 0.53 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END OR4X6

MACRO ACHCONX2
    CLASS CORE ;
    SIZE 5.2325 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN CON
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.8075 0.2295 4.688 0.272 ;
              RECT  4.2635 0.7175 4.628 0.76 ;
              RECT  4.2635 0.576 4.366 0.6325 ;
              RECT  4.3235 0.2295 4.366 0.6325 ;
              RECT  3.8995 0.7565 4.306 0.799 ;
              RECT  4.2635 0.576 4.306 0.799 ;
        END
    END CON
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0245 0.477 0.1445 0.767 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.117 0.491 1.2445 0.654 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.8115 0.548 5.137 0.6325 ;
        END
    END CI
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.2325 0.042 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.2325 1.209 ;
        END
    END VDD
END ACHCONX2

MACRO OAI21X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.502 0.8485 0.806 0.8905 ;
              RECT  0.7495 0.6925 0.806 0.8905 ;
              RECT  0.7495 0.304 0.7915 0.8905 ;
              RECT  0.647 0.304 0.7915 0.346 ;
              RECT  0.647 0.2615 0.689 0.346 ;
              RECT  0.502 0.8485 0.544 1.0465 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.424 0.537 0.4805 ;
              RECT  0.325 0.424 0.3815 0.622 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.7775 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OAI21X1

MACRO DLY3X4
    CLASS CORE ;
    SIZE 3.6765 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.424 1.23 0.516 ;
              RECT  1.117 0.431 1.1735 0.721 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.0575 0.3355 2.1425 0.378 ;
              RECT  2.0855 0.3355 2.128 0.912 ;
              RECT  1.739 0.424 2.128 0.4665 ;
              RECT  2.0575 0.3355 2.128 0.4665 ;
              RECT  1.796 0.424 1.838 0.912 ;
              RECT  1.739 0.3355 1.81 0.516 ;
              RECT  1.725 0.3355 1.81 0.378 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.6765 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.6765 0.042 ;
        END
    END VSS
END DLY3X4

MACRO TLATNSRX2
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8705 0.417 2.927 0.735 ;
              RECT  2.8175 0.3605 2.874 0.4735 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.3605 2.22 0.6925 ;
              RECT  2.146 0.636 2.2025 0.735 ;
        END
    END QN
    PIN GN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.012 0.5195 3.132 0.735 ;
              RECT  3.012 0.445 3.0685 0.735 ;
        END
    END GN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8805 0.53 1.937 0.8835 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.5585 1.3715 0.6505 ;
              RECT  1.0535 0.5585 1.3715 0.615 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5335 0.431 0.7245 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END TLATNSRX2

MACRO AND3XL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.286 0.806 0.979 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.6925 0.6645 0.7915 ;
              RECT  0.509 0.6925 0.6645 0.7495 ;
              RECT  0.509 0.537 0.5655 0.7495 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5585 0.325 0.643 ;
              RECT  0.2685 0.424 0.325 0.643 ;
              RECT  0.1835 0.5585 0.24 0.6925 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.424 0.0985 0.7775 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END AND3XL

MACRO DFFSXL
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.346 0.6645 0.721 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.159 0.3815 0.2155 0.721 ;
              RECT  0.042 0.424 0.2155 0.516 ;
        END
    END QN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.295 0.325 3.3515 0.6785 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.325 3.21 0.6785 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.576 1.545 0.6645 ;
              RECT  1.223 0.576 1.545 0.6325 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END DFFSXL

MACRO NAND4BBXL
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.788 0.2545 0.8305 0.979 ;
              RECT  0.4875 0.8695 0.8305 0.912 ;
              RECT  0.7495 0.6925 0.8305 0.912 ;
              RECT  0.392 0.2545 0.8305 0.2965 ;
              RECT  0.4875 0.8695 0.53 0.979 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.576 0.4945 0.799 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.4875 0.6645 0.6505 ;
              RECT  0.5655 0.5935 0.622 0.799 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0005 0.576 1.1065 0.781 ;
              RECT  0.9015 0.576 1.1065 0.6325 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.067 0.4415 0.1235 0.682 ;
              RECT  0.042 0.3535 0.0985 0.5265 ;
        END
    END BN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END NAND4BBXL

MACRO CLKBUFX16
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.902 0.403 1.9975 0.445 ;
              RECT  1.9335 0.6395 1.976 0.951 ;
              RECT  0.1625 0.4135 1.9335 0.456 ;
              RECT  0.1625 0.6395 1.976 0.682 ;
              RECT  1.6225 0.403 1.7075 0.456 ;
              RECT  1.644 0.6395 1.686 0.951 ;
              RECT  1.3325 0.403 1.4175 0.456 ;
              RECT  1.354 0.6395 1.3965 0.951 ;
              RECT  1.0425 0.403 1.1275 0.456 ;
              RECT  1.064 0.6395 1.1065 0.951 ;
              RECT  0.753 0.403 0.8375 0.456 ;
              RECT  0.774 0.6395 0.8165 0.951 ;
              RECT  0.463 0.403 0.548 0.456 ;
              RECT  0.484 0.6395 0.5265 0.951 ;
              RECT  0.1835 0.6395 0.24 0.7845 ;
              RECT  0.1835 0.6395 0.2365 0.951 ;
              RECT  0.194 0.371 0.2365 0.456 ;
              RECT  0.1625 0.4135 0.205 0.682 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.576 2.6585 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END CLKBUFX16

MACRO OAI221X1
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9225 0.7705 1.0605 0.813 ;
              RECT  1.018 0.2755 1.0605 0.813 ;
              RECT  0.8905 0.8485 0.965 1.0535 ;
              RECT  0.9225 0.7705 0.965 1.0535 ;
              RECT  0.5585 0.8485 0.965 0.8905 ;
              RECT  0.5585 0.8485 0.601 1.0465 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.7775 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.424 0.806 0.7775 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.332 0.9475 0.6855 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END OAI221X1

MACRO AND4XL
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.898 0.226 0.9475 0.88 ;
              RECT  0.8905 0.226 0.9475 0.3815 ;
              RECT  0.8305 0.226 0.9475 0.2685 ;
              RECT  0.8305 0.1835 0.873 0.2685 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.827 0.806 0.919 ;
              RECT  0.707 0.608 0.7635 0.8835 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4525 0.4525 0.523 0.6505 ;
              RECT  0.4525 0.4525 0.509 0.7915 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.311 0.4525 0.3815 0.6505 ;
              RECT  0.311 0.4525 0.3675 0.7915 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1555 0.4525 0.24 0.7775 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END AND4XL

MACRO OAI31X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.516 0.8485 0.806 0.8905 ;
              RECT  0.7635 0.2615 0.806 0.8905 ;
              RECT  0.7495 0.2615 0.806 0.3815 ;
              RECT  0.516 0.8485 0.5585 1.0465 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.1765 0.615 ;
              RECT  0.12 0.3745 0.1765 0.615 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.7775 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.424 0.523 0.7775 ;
        END
    END A2
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OAI31X1

MACRO OA21X1
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7635 0.403 0.919 0.445 ;
              RECT  0.7495 0.424 0.806 1.0285 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.3955 0.0985 0.7495 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.417 0.3815 0.7705 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.1555 0.523 0.509 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END OA21X1

MACRO DLY4X4
    CLASS CORE ;
    SIZE 4.384 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1645 0.5405 4.221 0.7495 ;
              RECT  4.1435 0.6925 4.2 0.873 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.735 0.6575 0.82 0.7 ;
              RECT  0.7565 0.346 0.799 0.7 ;
              RECT  0.4665 0.4735 0.799 0.516 ;
              RECT  0.4665 0.424 0.523 0.516 ;
              RECT  0.403 0.6575 0.509 0.7 ;
              RECT  0.4665 0.346 0.509 0.7 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.384 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.384 0.042 ;
        END
    END VSS
END DLY4X4

MACRO CLKXOR2X8
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.018 0.339 1.1135 0.3815 ;
              RECT  1.0535 0.647 1.096 0.9615 ;
              RECT  0.1835 0.647 1.096 0.689 ;
              RECT  0.18 0.35 1.05 0.392 ;
              RECT  0.7385 0.339 0.8235 0.392 ;
              RECT  0.7635 0.647 0.806 0.9615 ;
              RECT  0.449 0.339 0.5335 0.392 ;
              RECT  0.4735 0.647 0.516 0.9615 ;
              RECT  0.1835 0.35 0.24 0.516 ;
              RECT  0.1835 0.35 0.226 0.9615 ;
              RECT  0.18 0.3075 0.2225 0.392 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.5585 2.2485 0.615 ;
              RECT  2.1635 0.431 2.22 0.6505 ;
              RECT  1.923 0.431 2.22 0.4875 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3785 0.4415 1.435 0.714 ;
              RECT  1.2975 0.4415 1.435 0.5265 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END CLKXOR2X8

MACRO OR2X8
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.757 0.403 1.8525 0.445 ;
              RECT  0.951 0.4135 1.7885 0.456 ;
              RECT  1.7355 0.707 1.778 1.0215 ;
              RECT  0.866 0.707 1.778 0.7495 ;
              RECT  1.598 0.4135 1.6545 0.516 ;
              RECT  1.598 0.4135 1.64 0.7495 ;
              RECT  1.499 0.371 1.541 0.456 ;
              RECT  1.446 0.707 1.488 1.0215 ;
              RECT  1.1875 0.403 1.2725 0.456 ;
              RECT  1.156 0.707 1.1985 1.0215 ;
              RECT  0.898 0.403 0.9825 0.445 ;
              RECT  0.866 0.707 0.9085 1.0215 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.654 0.47 0.7105 ;
              RECT  0.325 0.654 0.3815 0.919 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.5265 0.682 0.583 ;
              RECT  0.1835 0.5585 0.2545 0.6505 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END OR2X8

MACRO DFFXL
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.7035 0.7455 0.788 ;
              RECT  0.6505 0.3675 0.707 0.4525 ;
              RECT  0.608 0.3955 0.6645 0.919 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1905 0.6645 0.247 0.7495 ;
              RECT  0.042 0.3815 0.247 0.4665 ;
              RECT  0.134 0.3815 0.1905 0.721 ;
              RECT  0.042 0.3815 0.1905 0.516 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7785 0.5975 2.9485 0.767 ;
              RECT  2.7785 0.5975 2.927 0.8375 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.919 0.576 1.1065 0.6325 ;
              RECT  0.919 0.438 0.9755 0.6325 ;
              RECT  0.8905 0.438 0.9755 0.5585 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END DFFXL

MACRO OAI2BB2X4
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.217 0.2155 3.302 0.258 ;
              RECT  2.563 0.2015 3.2525 0.2435 ;
              RECT  2.45 0.8165 3.1465 0.859 ;
              RECT  2.906 0.2015 2.991 0.258 ;
              RECT  2.5135 0.2155 2.5985 0.258 ;
              RECT  2.054 0.3285 2.556 0.371 ;
              RECT  2.5135 0.2155 2.556 0.371 ;
              RECT  1.7145 0.859 2.4925 0.9015 ;
              RECT  2.2025 0.3145 2.287 0.371 ;
              RECT  2.0045 0.8445 2.0965 0.9015 ;
              RECT  2.054 0.3285 2.0965 0.9015 ;
              RECT  1.7145 0.7845 1.9335 0.9015 ;
              RECT  1.7145 0.7845 1.757 0.9435 ;
              RECT  1.2055 0.7845 1.9335 0.827 ;
              RECT  1.2055 0.7845 1.248 0.8695 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.181 0.4415 2.5065 0.4985 ;
              RECT  2.3225 0.4415 2.379 0.5265 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.164 0.59 3.3125 0.6325 ;
              RECT  2.167 0.5975 3.2065 0.6395 ;
              RECT  2.2095 0.5975 2.379 0.767 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.484 0.3815 0.8375 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.484 0.24 0.8375 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END OAI2BB2X4

MACRO EDFFX1
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.7335 0.3815 3.7755 0.912 ;
              RECT  3.719 0.424 3.7755 0.516 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.3815 3.21 0.912 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8705 0.689 2.927 0.7845 ;
              RECT  2.287 0.7635 2.913 0.806 ;
              RECT  2.0965 1.0285 2.3295 1.071 ;
              RECT  2.287 0.491 2.3295 1.071 ;
              RECT  2.245 0.491 2.3295 0.5335 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.5135 0.569 2.8 0.6255 ;
              RECT  2.5135 0.569 2.662 0.6925 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.3815 0.7845 ;
              RECT  0.212 0.6925 0.3815 0.7495 ;
              RECT  0.212 0.544 0.2685 0.7495 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END EDFFX1

MACRO HOLDX1
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.615 0.3815 0.6645 0.721 ;
              RECT  0.24 0.6505 0.6645 0.6925 ;
              RECT  0.608 0.5585 0.6645 0.6925 ;
              RECT  0.24 0.523 0.2825 0.6925 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END HOLDX1

MACRO TLATNTSCAX8
    CLASS CORE ;
    SIZE 3.6765 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4715 0.3535 3.514 0.993 ;
              RECT  2.588 0.6785 3.514 0.721 ;
              RECT  2.9235 0.3955 3.514 0.438 ;
              RECT  3.1605 0.385 3.2455 0.438 ;
              RECT  3.1815 0.6785 3.224 0.993 ;
              RECT  2.8705 0.385 2.9555 0.4275 ;
              RECT  2.892 0.6785 2.934 0.993 ;
              RECT  2.602 0.364 2.6445 0.993 ;
              RECT  2.588 0.6785 2.6445 0.7845 ;
        END
    END ECK
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.477 0.424 0.5335 0.661 ;
              RECT  0.4665 0.318 0.523 0.516 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3145 0.318 0.3815 0.516 ;
              RECT  0.3145 0.318 0.371 0.661 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0455 0.3285 0.1305 0.6325 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.6765 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.6765 0.042 ;
        END
    END VSS
END TLATNTSCAX8

MACRO ANTENNA
    CLASS CORE ;
    SIZE 0.424 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.424 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.424 0.042 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.2755 0.24 0.898 ;
        END
    END A
END ANTENNA

MACRO OAI2BB2X1
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0145 0.8445 1.4845 0.887 ;
              RECT  1.442 0.311 1.4845 0.887 ;
              RECT  1.4105 0.2685 1.453 0.3535 ;
              RECT  1.2335 0.8445 1.276 0.9295 ;
              RECT  1.0145 0.8445 1.276 0.9015 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5555 0.5335 1.6545 0.6395 ;
              RECT  1.598 0.3285 1.6545 0.6395 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.4205 1.3715 0.774 ;
        END
    END B1
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4415 0.7105 0.647 0.781 ;
              RECT  0.4415 0.576 0.502 0.781 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3145 0.576 0.371 0.781 ;
              RECT  0.166 0.576 0.371 0.6325 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END OAI2BB2X1

MACRO CLKINVX1
    CLASS CORE ;
    SIZE 0.424 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.3605 0.24 0.912 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.417 0.113 0.7565 ;
              RECT  0.042 0.417 0.113 0.5585 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.424 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.424 0.042 ;
        END
    END VSS
END CLKINVX1

MACRO SDFFHQX2
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.212 0.3815 0.2545 0.9435 ;
              RECT  0.1835 0.5585 0.2545 0.6505 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.56 0.576 3.652 0.6325 ;
              RECT  3.5955 0.3535 3.638 0.6325 ;
              RECT  2.966 0.3535 3.638 0.3955 ;
              RECT  3.553 0.576 3.652 0.6185 ;
              RECT  3.1395 0.3535 3.224 0.4735 ;
              RECT  2.966 0.3535 3.0085 0.622 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.295 0.555 3.4825 0.689 ;
              RECT  3.4255 0.4665 3.4825 0.689 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7255 0.456 2.782 0.569 ;
              RECT  2.588 0.456 2.782 0.516 ;
              RECT  2.588 0.3535 2.6445 0.516 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6645 0.576 0.721 ;
              RECT  0.449 0.629 0.576 0.721 ;
              RECT  0.325 0.6645 0.3815 0.788 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END SDFFHQX2

MACRO SDFFSRHQX8
    CLASS CORE ;
    SIZE 6.788 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  6.5475 0.424 6.604 0.516 ;
              RECT  5.9395 0.424 6.604 0.4665 ;
              RECT  5.9395 0.424 5.982 0.622 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  6.208 0.5795 6.477 0.6785 ;
              RECT  6.247 0.537 6.477 0.6785 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.699 0.3145 5.7555 0.668 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.572 0.4415 5.6285 0.622 ;
              RECT  5.3985 0.4415 5.6285 0.4985 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.705 0.905 4.2425 0.9475 ;
              RECT  3.705 0.8025 3.7475 0.9475 ;
              RECT  3.4365 0.8025 3.7475 0.8445 ;
              RECT  2.8705 0.9225 3.4785 0.965 ;
              RECT  3.4365 0.8025 3.4785 0.965 ;
              RECT  2.8705 0.675 2.913 0.965 ;
              RECT  2.206 0.675 2.913 0.7175 ;
              RECT  2.206 0.576 2.2485 0.7175 ;
              RECT  2.1635 0.5585 2.22 0.6505 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8135 0.5585 2.093 0.615 ;
              RECT  1.8135 0.5585 1.955 0.689 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.926 0.636 0.9685 0.951 ;
              RECT  0.926 0.3745 0.9685 0.4595 ;
              RECT  0.894 0.417 0.9365 0.6785 ;
              RECT  0.636 0.523 0.9365 0.5655 ;
              RECT  0.636 0.3815 0.6785 0.951 ;
              RECT  0.042 0.424 0.6785 0.4665 ;
              RECT  0.346 0.3815 0.3885 0.951 ;
              RECT  0.0565 0.3815 0.0985 0.951 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.788 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.788 0.042 ;
        END
    END VSS
END SDFFSRHQX8

MACRO CLKXOR2X2
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.265 0.8165 0.3075 0.9015 ;
              RECT  0.1975 0.35 0.3075 0.392 ;
              RECT  0.265 0.3075 0.3075 0.392 ;
              RECT  0.1975 0.8165 0.3075 0.859 ;
              RECT  0.1975 0.35 0.24 0.859 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9435 0.576 1.262 0.6185 ;
              RECT  1.0145 0.576 1.1065 0.6325 ;
              RECT  0.7495 0.583 1.1065 0.6255 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.509 0.576 0.5655 0.8445 ;
              RECT  0.424 0.576 0.5655 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END CLKXOR2X2

MACRO OAI221X4
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.998 0.5585 3.0685 0.6505 ;
              RECT  2.9165 0.7565 3.0405 0.799 ;
              RECT  2.998 0.378 3.0405 0.799 ;
              RECT  2.6905 0.4345 3.0405 0.477 ;
              RECT  2.98 0.378 3.0405 0.477 ;
              RECT  2.9165 0.7565 2.959 1.032 ;
              RECT  0.403 0.8555 2.959 0.898 ;
              RECT  2.6905 0.378 2.7325 0.477 ;
              RECT  2.6265 0.7565 2.669 1.032 ;
              RECT  2.153 0.8555 2.1955 0.94 ;
              RECT  1.7145 0.8555 1.757 0.94 ;
              RECT  1.025 0.8555 1.0675 0.94 ;
              RECT  0.403 0.8555 0.445 0.94 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.7035 1.2405 0.7455 ;
              RECT  1.1985 0.643 1.2405 0.7455 ;
              RECT  0.714 0.661 0.7565 0.7455 ;
              RECT  0.1975 0.5585 0.24 0.7455 ;
              RECT  0.1555 0.608 0.24 0.6505 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4775 0.742 2.503 0.7845 ;
              RECT  2.4465 0.643 2.503 0.7845 ;
              RECT  1.9585 0.6645 2.0435 0.7845 ;
              RECT  1.4775 0.6185 1.52 0.7845 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4345 0.548 1.0425 0.59 ;
              RECT  0.4345 0.548 0.5405 0.6325 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.146 0.576 2.2375 0.6325 ;
              RECT  1.7465 0.548 2.206 0.59 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.5735 0.576 2.927 0.6325 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END OAI221X4

MACRO XNOR3X1
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.287 0.576 2.379 0.661 ;
              RECT  2.287 0.47 2.3295 0.661 ;
              RECT  2.068 0.47 2.3295 0.5125 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.4735 0.3815 0.7455 ;
              RECT  0.2895 0.4275 0.346 0.53 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.4345 0.106 0.781 ;
              RECT  0.042 0.5585 0.106 0.6505 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.998 0.6575 3.0865 0.7 ;
              RECT  3.044 0.3075 3.0865 0.7 ;
              RECT  2.9945 0.3075 3.0865 0.364 ;
        END
    END Y
END XNOR3X1

MACRO SEDFFXL
    CLASS CORE ;
    SIZE 5.091 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.729 0.7635 2.814 0.82 ;
              RECT  2.729 0.2965 2.786 0.82 ;
              RECT  2.7185 0.265 2.775 0.3535 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1985 0.4595 1.255 0.8555 ;
              RECT  1.1525 0.424 1.23 0.4805 ;
              RECT  1.1525 0.339 1.209 0.4805 ;
              RECT  1.1735 0.4595 1.255 0.516 ;
        END
    END QN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.8505 0.5585 5.0695 0.643 ;
              RECT  4.8505 0.5585 4.907 0.7495 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4465 0.403 2.503 0.7565 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.576 1.7815 0.6325 ;
              RECT  1.725 0.5195 1.7815 0.6325 ;
              RECT  1.598 0.5195 1.6545 0.689 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.569 0.4985 0.675 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9085 0.2295 0.951 0.6575 ;
              RECT  0.4985 0.2295 0.951 0.272 ;
              RECT  0.569 0.456 0.6115 0.544 ;
              RECT  0.194 0.456 0.6115 0.4985 ;
              RECT  0.449 0.4415 0.5405 0.4985 ;
              RECT  0.4985 0.2295 0.5405 0.4985 ;
              RECT  0.194 0.456 0.2365 0.544 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.091 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.091 0.042 ;
        END
    END VSS
END SEDFFXL

MACRO OA22X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0465 0.371 1.1415 0.4135 ;
              RECT  1.0465 0.371 1.0885 0.516 ;
              RECT  1.018 0.4735 1.0605 0.94 ;
              RECT  1.032 0.424 1.0885 0.516 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.6925 0.9475 0.7845 ;
              RECT  0.707 0.6925 0.9475 0.7495 ;
              RECT  0.707 0.615 0.7635 0.7495 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.24 0.7845 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.4525 0.523 0.806 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OA22X1

MACRO AOI211X1
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7315 0.7915 0.919 0.834 ;
              RECT  0.8765 0.339 0.919 0.834 ;
              RECT  0.445 0.339 0.919 0.3815 ;
              RECT  0.7495 0.2895 0.806 0.3815 ;
              RECT  0.7315 0.7915 0.774 1.0465 ;
              RECT  0.41 0.311 0.4945 0.3535 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.424 0.3815 0.7775 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.4525 0.5935 0.509 ;
              RECT  0.4665 0.4525 0.523 0.735 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.5585 0.806 0.721 ;
              RECT  0.6645 0.5585 0.806 0.615 ;
              RECT  0.6645 0.4525 0.721 0.615 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END AOI211X1

MACRO TLATX4
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.711 0.371 2.0855 0.4135 ;
              RECT  2.0435 0.3285 2.0855 0.4135 ;
              RECT  1.916 0.7245 1.9585 0.958 ;
              RECT  1.598 0.7245 1.9585 0.767 ;
              RECT  1.598 0.6925 1.7535 0.767 ;
              RECT  1.711 0.3285 1.7535 0.767 ;
              RECT  1.598 0.6925 1.6685 0.958 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7565 0.682 0.799 0.958 ;
              RECT  0.3815 0.371 0.7565 0.4135 ;
              RECT  0.714 0.3285 0.7565 0.4135 ;
              RECT  0.4665 0.682 0.799 0.7245 ;
              RECT  0.4805 0.371 0.523 0.7245 ;
              RECT  0.4665 0.5585 0.509 0.958 ;
              RECT  0.3815 0.3285 0.424 0.4135 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.5585 3.21 0.753 ;
              RECT  2.9945 0.5585 3.21 0.6505 ;
        END
    END D
    PIN G
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.325 0.24 0.6785 ;
        END
    END G
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END TLATX4

MACRO BUFX20
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3685 0.647 2.411 0.9615 ;
              RECT  0.042 0.4205 2.411 0.463 ;
              RECT  2.3685 0.251 2.411 0.463 ;
              RECT  0.042 0.647 2.411 0.689 ;
              RECT  2.0785 0.647 2.121 0.9615 ;
              RECT  2.0785 0.251 2.121 0.463 ;
              RECT  1.7885 0.647 1.831 0.9615 ;
              RECT  1.7885 0.251 1.831 0.463 ;
              RECT  1.499 0.647 1.541 0.9615 ;
              RECT  1.499 0.251 1.541 0.463 ;
              RECT  1.209 0.647 1.2515 0.9615 ;
              RECT  1.209 0.251 1.2515 0.463 ;
              RECT  0.919 0.647 0.9615 0.9615 ;
              RECT  0.919 0.251 0.9615 0.463 ;
              RECT  0.629 0.647 0.6715 0.9615 ;
              RECT  0.629 0.251 0.6715 0.463 ;
              RECT  0.339 0.647 0.3815 0.9615 ;
              RECT  0.339 0.251 0.3815 0.463 ;
              RECT  0.042 0.4205 0.0985 0.689 ;
              RECT  0.042 0.251 0.0915 0.9615 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.74 0.576 3.0935 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END BUFX20

MACRO XNOR2XL
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.424 0.2085 0.4805 ;
              RECT  0.152 0.3425 0.2085 0.4805 ;
              RECT  0.0845 0.424 0.141 0.7775 ;
              RECT  0.042 0.424 0.141 0.516 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.898 0.576 1.2515 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.456 0.615 ;
              RECT  0.3995 0.4805 0.456 0.615 ;
              RECT  0.325 0.5585 0.3815 0.76 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END XNOR2XL

MACRO OR4X1
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.2895 0.9475 0.3815 ;
              RECT  0.8765 0.279 0.919 0.979 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3605 0.4665 0.417 0.7565 ;
              RECT  0.325 0.6925 0.3815 0.7845 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.233 0.417 0.2895 0.615 ;
              RECT  0.1835 0.5585 0.24 0.721 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.417 0.113 0.562 ;
              RECT  0.021 0.5195 0.0845 0.735 ;
        END
    END D
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.601 0.484 0.806 0.5405 ;
              RECT  0.7495 0.3355 0.806 0.5405 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END OR4X1

MACRO OAI211XL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.841 0.806 0.9755 ;
              RECT  0.735 0.2085 0.7775 0.926 ;
              RECT  0.41 0.8835 0.806 0.926 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5655 0.24 0.919 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.4595 0.3815 0.813 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.47 0.463 0.5265 0.813 ;
              RECT  0.4665 0.463 0.5265 0.6505 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.7775 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OAI211XL

MACRO BUFX4
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4735 0.2825 0.5585 0.325 ;
              RECT  0.4945 0.6925 0.537 0.9685 ;
              RECT  0.1625 0.2965 0.509 0.339 ;
              RECT  0.1625 0.6925 0.537 0.735 ;
              RECT  0.1835 0.6925 0.24 0.7845 ;
              RECT  0.1835 0.6925 0.2365 0.9685 ;
              RECT  0.194 0.2545 0.2365 0.339 ;
              RECT  0.1625 0.2965 0.205 0.735 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.5515 0.728 0.608 ;
              RECT  0.6715 0.523 0.728 0.608 ;
              RECT  0.608 0.5515 0.6645 0.813 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END BUFX4

MACRO CLKINVX4
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.6925 0.6645 0.7845 ;
              RECT  0.608 0.438 0.6505 0.7845 ;
              RECT  0.5725 0.7035 0.615 0.9435 ;
              RECT  0.2825 0.438 0.6505 0.4805 ;
              RECT  0.5725 0.3815 0.615 0.4805 ;
              RECT  0.2825 0.7035 0.6645 0.7455 ;
              RECT  0.2825 0.7035 0.325 0.9435 ;
              RECT  0.2825 0.3815 0.325 0.4805 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.576 0.537 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END CLKINVX4

MACRO AOI33X4
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5495 0.767 3.592 0.852 ;
              RECT  2.39 0.767 3.592 0.8095 ;
              RECT  3.2595 0.767 3.302 0.852 ;
              RECT  0.675 0.2365 3.2525 0.279 ;
              RECT  2.9695 0.767 3.012 0.852 ;
              RECT  2.6795 0.767 2.722 0.852 ;
              RECT  2.39 0.7035 2.432 0.852 ;
              RECT  2.1 0.7035 2.432 0.7455 ;
              RECT  2.1 0.576 2.1425 0.788 ;
              RECT  1.8665 0.576 2.1425 0.6325 ;
              RECT  1.8665 0.5585 1.937 0.6505 ;
              RECT  1.8665 0.2365 1.909 0.6505 ;
        END
    END Y
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.576 1.5305 0.6325 ;
              RECT  1.4385 0.576 1.5025 0.661 ;
              RECT  0.8695 0.654 1.481 0.6965 ;
              RECT  0.8695 0.5975 0.912 0.6965 ;
              RECT  0.689 0.5975 0.912 0.6395 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.026 0.59 3.231 0.6325 ;
              RECT  2.503 0.654 3.0685 0.6965 ;
              RECT  3.026 0.59 3.0685 0.6965 ;
              RECT  2.503 0.576 2.5455 0.6965 ;
              RECT  2.4285 0.576 2.5455 0.6325 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4365 0.548 3.5 0.6325 ;
              RECT  3.4365 0.548 3.493 0.6505 ;
              RECT  3.302 0.548 3.5 0.59 ;
              RECT  3.302 0.477 3.3445 0.59 ;
              RECT  2.913 0.477 3.3445 0.5195 ;
              RECT  2.616 0.5405 2.9555 0.583 ;
              RECT  2.913 0.477 2.9555 0.583 ;
              RECT  2.616 0.463 2.6585 0.583 ;
              RECT  2.1705 0.463 2.6585 0.5055 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3255 0.463 1.6685 0.5055 ;
              RECT  0.9825 0.5405 1.368 0.583 ;
              RECT  1.3255 0.463 1.368 0.583 ;
              RECT  0.9825 0.484 1.025 0.583 ;
              RECT  0.4805 0.484 1.025 0.5265 ;
              RECT  0.4665 0.5585 0.523 0.6505 ;
              RECT  0.4805 0.484 0.523 0.6505 ;
              RECT  0.424 0.5585 0.523 0.601 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.35 1.796 0.516 ;
              RECT  0.311 0.35 1.796 0.392 ;
              RECT  1.096 0.35 1.1805 0.47 ;
              RECT  0.311 0.35 0.3535 0.491 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5705 0.35 3.613 0.4985 ;
              RECT  2.054 0.35 3.613 0.392 ;
              RECT  2.7575 0.35 2.8425 0.47 ;
              RECT  1.9795 0.4135 2.0965 0.47 ;
              RECT  2.054 0.35 2.0965 0.47 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END AOI33X4

MACRO TBUFX16
    CLASS CORE ;
    SIZE 6.3635 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.9995 0.728 6.042 1.004 ;
              RECT  4.002 0.728 6.042 0.7705 ;
              RECT  5.918 0.2615 5.9605 0.7705 ;
              RECT  5.3385 0.318 5.9605 0.3605 ;
              RECT  5.7095 0.728 5.752 1.004 ;
              RECT  5.6285 0.2615 5.6705 0.3605 ;
              RECT  5.4195 0.728 5.462 1.004 ;
              RECT  5.3385 0.2615 5.381 0.3605 ;
              RECT  5.13 0.728 5.172 1.004 ;
              RECT  5.0485 0.2615 5.091 0.7705 ;
              RECT  4.7585 0.318 5.091 0.3605 ;
              RECT  4.84 0.728 4.8825 1.004 ;
              RECT  4.7585 0.2615 4.801 0.3605 ;
              RECT  4.55 0.728 4.5925 1.004 ;
              RECT  4.179 0.318 4.511 0.3605 ;
              RECT  4.4685 0.2615 4.511 0.3605 ;
              RECT  4.26 0.318 4.3025 1.004 ;
              RECT  4.179 0.2615 4.221 0.3605 ;
              RECT  4.002 0.5585 4.0585 0.7705 ;
              RECT  4.002 0.318 4.0445 0.795 ;
              RECT  3.97 0.753 4.0125 1.004 ;
              RECT  3.889 0.318 4.0445 0.3605 ;
              RECT  3.889 0.2615 3.9315 0.3605 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4785 0.449 3.6625 0.491 ;
              RECT  2.1635 0.431 3.521 0.4735 ;
              RECT  2.1635 0.318 2.206 0.4735 ;
              RECT  1.8135 0.2895 2.1775 0.332 ;
              RECT  2.135 0.318 2.206 0.3605 ;
              RECT  1.587 0.477 1.856 0.5195 ;
              RECT  1.8135 0.2895 1.856 0.5195 ;
              RECT  1.6545 0.477 1.697 0.5975 ;
              RECT  1.587 0.2895 1.6295 0.5195 ;
              RECT  1.276 0.2895 1.6295 0.332 ;
              RECT  1.0075 0.456 1.3185 0.4985 ;
              RECT  1.276 0.2895 1.3185 0.4985 ;
              RECT  1.1275 0.456 1.17 0.5865 ;
              RECT  1.0075 0.2895 1.05 0.4985 ;
              RECT  0.7315 0.2895 1.05 0.332 ;
              RECT  0.7315 0.576 0.8235 0.6325 ;
              RECT  0.4985 0.6575 0.774 0.7 ;
              RECT  0.7315 0.2895 0.774 0.7 ;
              RECT  0.364 0.615 0.5405 0.6575 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6185 0.502 0.661 0.5865 ;
              RECT  0.1835 0.502 0.661 0.544 ;
              RECT  0.1835 0.502 0.293 0.6505 ;
        END
    END OE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.3635 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.3635 0.042 ;
        END
    END VSS
END TBUFX16

MACRO SDFFRX1
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.622 0.3815 0.6645 0.94 ;
              RECT  0.608 0.424 0.6645 0.516 ;
              RECT  0.6115 0.3815 0.6645 0.516 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.148 0.3815 0.205 0.912 ;
              RECT  0.042 0.424 0.205 0.516 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.285 0.424 4.3415 0.516 ;
              RECT  4.285 0.3285 4.327 0.516 ;
              RECT  3.8215 0.3285 4.327 0.371 ;
              RECT  3.6345 0.477 3.864 0.5195 ;
              RECT  3.8215 0.3285 3.864 0.5195 ;
              RECT  3.6345 0.477 3.6765 0.562 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.935 0.4415 4.214 0.5265 ;
              RECT  3.935 0.4415 3.9915 0.5725 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.295 0.35 3.4505 0.4065 ;
              RECT  3.295 0.35 3.3515 0.6045 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2725 0.5195 1.5235 0.576 ;
              RECT  1.2725 0.5195 1.389 0.6785 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6925 0.905 0.7845 ;
              RECT  0.8485 0.53 0.905 0.7845 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END SDFFRX1

MACRO DFFSRHQX8
    CLASS CORE ;
    SIZE 5.515 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.275 0.463 5.3315 0.8165 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.833 0.35 4.932 0.4985 ;
              RECT  4.7835 0.4415 4.868 0.6115 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.7335 0.9755 3.9525 1.018 ;
              RECT  3.7335 0.8625 3.7755 1.018 ;
              RECT  3.4645 0.8625 3.7755 0.905 ;
              RECT  2.7575 0.9085 3.507 0.951 ;
              RECT  3.4645 0.8625 3.507 0.951 ;
              RECT  2.7575 0.795 2.8 0.951 ;
              RECT  2.418 0.795 2.8 0.8375 ;
              RECT  2.1775 0.852 2.4605 0.894 ;
              RECT  2.418 0.795 2.4605 0.894 ;
              RECT  2.1775 0.5585 2.22 0.894 ;
              RECT  2.1635 0.5585 2.22 0.6505 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8805 0.424 1.937 0.7775 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.926 0.636 0.9685 0.951 ;
              RECT  0.926 0.3745 0.9685 0.4595 ;
              RECT  0.894 0.417 0.9365 0.6785 ;
              RECT  0.636 0.523 0.9365 0.5655 ;
              RECT  0.636 0.3815 0.6785 0.951 ;
              RECT  0.042 0.456 0.6785 0.4985 ;
              RECT  0.346 0.3815 0.3885 0.951 ;
              RECT  0.0565 0.3815 0.0985 0.951 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.515 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.515 0.042 ;
        END
    END VSS
END DFFSRHQX8

MACRO AOI222X2
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.015 0.7175 2.0575 0.8025 ;
              RECT  1.725 0.721 2.0575 0.7635 ;
              RECT  0.4985 0.318 1.8915 0.3605 ;
              RECT  1.725 0.7105 1.7675 0.8165 ;
              RECT  0.905 0.7105 1.7675 0.753 ;
              RECT  0.905 0.318 0.9475 0.753 ;
              RECT  0.8905 0.5585 0.9475 0.6505 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.576 1.5095 0.6325 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5585 0.59 0.6505 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8065 0.576 1.937 0.6325 ;
              RECT  1.8065 0.5585 1.9265 0.6505 ;
        END
    END C1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6115 0.449 0.7495 0.5055 ;
              RECT  0.357 0.431 0.6715 0.4875 ;
              RECT  0.166 0.4415 0.3955 0.523 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.064 0.449 1.5095 0.5055 ;
              RECT  1.2975 0.4415 1.389 0.5055 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.008 0.4805 2.1315 0.523 ;
              RECT  1.58 0.4415 2.0505 0.484 ;
              RECT  1.58 0.4415 1.697 0.5055 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END AOI222X2

MACRO NAND2BX1
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.7105 0.106 0.767 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.417 0.569 0.544 0.682 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.438 0.1165 0.4985 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.5655 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.5655 0.042 ;
        END
    END VSS
END NAND2BX1

MACRO AOI211X4
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4005 0.7385 2.443 0.9015 ;
              RECT  2.3295 0.3145 2.4145 0.357 ;
              RECT  2.1105 0.7385 2.443 0.781 ;
              RECT  0.5865 0.3285 2.365 0.371 ;
              RECT  2.1105 0.7035 2.153 0.9015 ;
              RECT  1.347 0.7035 2.153 0.7455 ;
              RECT  2.0185 0.3145 2.1035 0.371 ;
              RECT  1.7075 0.3145 1.7925 0.371 ;
              RECT  1.368 0.3145 1.453 0.371 ;
              RECT  1.347 0.3285 1.389 0.7455 ;
              RECT  1.2975 0.4415 1.389 0.4985 ;
              RECT  0.9755 0.3145 1.0605 0.371 ;
              RECT  0.537 0.3145 0.622 0.357 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.576 1.0075 0.6325 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.46 0.576 1.8135 0.6325 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3225 0.4415 2.379 0.583 ;
              RECT  2.1105 0.4415 2.379 0.4985 ;
        END
    END C0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1625 0.456 1.2265 0.4985 ;
              RECT  0.166 0.4415 0.258 0.4985 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END AOI211X4

MACRO BMXIX4
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN M1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.283 0.562 1.7005 0.6045 ;
              RECT  1.658 0.5195 1.7005 0.6045 ;
              RECT  1.283 0.4415 1.389 0.6045 ;
              RECT  1.283 0.134 1.3255 0.6045 ;
              RECT  1.124 0.134 1.3255 0.1765 ;
              RECT  1.0815 0.0915 1.1665 0.134 ;
        END
    END M1
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.318 0.9475 0.6715 ;
        END
    END A
    PIN S
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.9015 1.474 0.9435 ;
              RECT  0.7495 0.8555 0.7915 0.9435 ;
              RECT  0.4665 0.8555 0.7915 0.898 ;
              RECT  0.4665 0.6925 0.523 0.898 ;
              RECT  0.4665 0.537 0.509 0.898 ;
              RECT  0.2825 0.537 0.509 0.5795 ;
        END
    END S
    PIN M0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3535 0.9685 0.6785 1.011 ;
              RECT  0.3535 0.859 0.3955 1.011 ;
              RECT  0.166 0.859 0.3955 0.9015 ;
              RECT  0.166 0.8445 0.258 0.9015 ;
              RECT  0.166 0.5405 0.2085 0.9015 ;
        END
    END M0
    PIN PPN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.2985 0.3815 3.341 0.912 ;
              RECT  3.0085 0.4735 3.341 0.516 ;
              RECT  3.0085 0.424 3.0685 0.516 ;
              RECT  3.0085 0.3815 3.051 0.912 ;
        END
    END PPN
    PIN X2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4285 0.979 2.5205 1.0355 ;
              RECT  2.2375 0.979 2.5205 1.0215 ;
              RECT  2.2375 0.5195 2.28 1.0215 ;
              RECT  2.174 0.5195 2.28 0.6045 ;
        END
    END X2
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END BMXIX4

MACRO MX4XL
    CLASS CORE ;
    SIZE 2.9695 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0845 0.2895 0.141 0.3745 ;
              RECT  0.042 0.5585 0.113 0.721 ;
              RECT  0.042 0.318 0.0985 0.721 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.478 0.583 2.8035 0.6325 ;
              RECT  2.687 0.576 2.8035 0.6325 ;
              RECT  2.478 0.583 2.5205 1.018 ;
              RECT  1.824 0.9755 2.5205 1.018 ;
              RECT  2.4355 0.583 2.8035 0.6255 ;
              RECT  1.6475 1.011 1.8665 1.0535 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.45 0.4415 2.8035 0.4985 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.04 0.555 2.0965 0.7915 ;
              RECT  1.923 0.555 2.0965 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.796 0.7105 1.969 0.767 ;
              RECT  1.796 0.5585 1.8525 0.767 ;
              RECT  1.7675 0.5585 1.8525 0.615 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.4735 1.3715 0.827 ;
        END
    END D
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5585 0.3815 0.615 ;
              RECT  0.325 0.438 0.3815 0.615 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END S1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.9695 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.9695 0.042 ;
        END
    END VSS
END MX4XL

MACRO TLATX2
    CLASS CORE ;
    SIZE 2.5455 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.5455 0.042 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.5455 1.209 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2545 0.5195 0.417 0.576 ;
              RECT  0.2545 0.5195 0.3995 0.767 ;
        END
    END D
    PIN G
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2975 0.576 1.4245 0.767 ;
        END
    END G
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.2895 1.6545 0.3815 ;
              RECT  1.598 0.2895 1.64 0.9225 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.325 2.3615 0.9225 ;
        END
    END Q
END TLATX2

MACRO TBUFX8
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.623 0.3745 3.2455 0.417 ;
              RECT  3.203 0.318 3.2455 0.417 ;
              RECT  3.1675 0.3745 3.21 0.912 ;
              RECT  2.4465 0.636 3.21 0.6785 ;
              RECT  2.913 0.318 2.9555 0.417 ;
              RECT  2.8775 0.636 2.92 0.912 ;
              RECT  2.623 0.318 2.6655 0.417 ;
              RECT  2.588 0.636 2.63 0.912 ;
              RECT  2.4465 0.5585 2.503 0.6785 ;
              RECT  2.298 0.7 2.489 0.742 ;
              RECT  2.4465 0.41 2.489 0.742 ;
              RECT  2.333 0.41 2.489 0.4525 ;
              RECT  2.333 0.318 2.3755 0.4525 ;
              RECT  2.298 0.7 2.3405 0.912 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.001 0.187 2.1425 0.2295 ;
              RECT  0.94 0.1905 2.0435 0.233 ;
              RECT  0.417 0.608 0.9825 0.6505 ;
              RECT  0.94 0.1905 0.9825 0.6505 ;
              RECT  0.449 0.576 0.5405 0.6505 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.827 0.4525 0.8695 0.537 ;
              RECT  0.1835 0.463 0.8695 0.5055 ;
              RECT  0.6115 0.463 0.6965 0.5335 ;
              RECT  0.1555 0.608 0.24 0.6505 ;
              RECT  0.1835 0.463 0.24 0.6505 ;
        END
    END OE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END TBUFX8

MACRO NAND2BX4
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0455 0.385 0.1025 0.4415 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.272 0.654 0.3285 0.7105 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3115 0.555 1.368 0.6575 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END NAND2BX4

MACRO SDFFQXL
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.2895 0.0985 0.9545 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9945 0.4415 3.0865 0.4985 ;
              RECT  2.662 0.4415 3.0865 0.484 ;
              RECT  2.6195 0.6395 2.7045 0.682 ;
              RECT  2.662 0.4415 2.7045 0.682 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.775 0.608 3.09 0.6645 ;
              RECT  2.775 0.569 2.945 0.6645 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.082 0.576 2.4355 0.6325 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.233 0.562 0.2895 0.7495 ;
              RECT  0.1835 0.6925 0.24 0.866 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END SDFFQXL

MACRO AOI33X2
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.831 0.7385 1.8735 0.8235 ;
              RECT  1.2265 0.7385 1.8735 0.781 ;
              RECT  1.527 0.7385 1.5695 0.8235 ;
              RECT  0.5335 0.2365 1.552 0.279 ;
              RECT  1.2265 0.7245 1.269 0.8235 ;
              RECT  1.0145 0.7245 1.269 0.767 ;
              RECT  1.0145 0.7105 1.1065 0.767 ;
              RECT  1.0605 0.2365 1.103 0.767 ;
        END
    END Y
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.576 0.82 0.6325 ;
              RECT  0.484 0.576 0.682 0.6505 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3395 0.576 1.6685 0.6325 ;
              RECT  1.3395 0.576 1.513 0.6575 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.463 1.796 0.6505 ;
              RECT  1.301 0.463 1.796 0.5055 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2965 0.463 0.7845 0.5055 ;
              RECT  0.325 0.463 0.3815 0.6505 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.424 0.9475 0.5195 ;
              RECT  0.8905 0.35 0.933 0.5195 ;
              RECT  0.1835 0.35 0.933 0.392 ;
              RECT  0.1835 0.35 0.226 0.5125 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8665 0.35 1.909 0.5195 ;
              RECT  1.1875 0.35 1.909 0.392 ;
              RECT  1.1735 0.424 1.23 0.5195 ;
              RECT  1.1875 0.35 1.23 0.5195 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END AOI33X2

MACRO ADDFX1
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.729 0.2895 2.786 0.3815 ;
              RECT  2.729 0.2895 2.7715 0.7495 ;
              RECT  2.687 0.707 2.729 0.9825 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2435 0.636 0.286 0.912 ;
              RECT  0.0565 0.41 0.286 0.4525 ;
              RECT  0.2435 0.3535 0.286 0.4525 ;
              RECT  0.042 0.636 0.286 0.6785 ;
              RECT  0.042 0.5585 0.0985 0.6785 ;
              RECT  0.0565 0.41 0.0985 0.6785 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.5795 2.3755 0.622 ;
              RECT  0.788 0.6115 1.481 0.654 ;
              RECT  1.2975 0.6115 1.389 0.767 ;
              RECT  0.788 0.569 0.8305 0.654 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4465 0.4665 2.503 0.6505 ;
              RECT  1.3505 0.4665 2.503 0.509 ;
              RECT  0.9015 0.477 1.393 0.5195 ;
              RECT  0.6715 0.456 0.9435 0.4985 ;
              RECT  0.629 0.4735 0.714 0.516 ;
        END
    END A
    PIN CI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1275 0.3535 2.2485 0.3955 ;
              RECT  1.1275 0.3075 1.248 0.3955 ;
              RECT  1.1275 0.3075 1.17 0.4065 ;
        END
    END CI
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END ADDFX1

MACRO SDFFHQX8
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.483 0.4415 4.525 0.5265 ;
              RECT  4.4085 0.4415 4.525 0.4985 ;
              RECT  3.977 0.456 4.525 0.4985 ;
              RECT  3.9135 0.491 4.0195 0.5335 ;
              RECT  3.9135 0.491 3.956 0.682 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.147 0.569 4.412 0.6255 ;
              RECT  4.147 0.569 4.359 0.714 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.673 0.5585 3.7295 0.7175 ;
              RECT  3.5775 0.5585 3.7295 0.6505 ;
              RECT  3.5775 0.4595 3.6345 0.6505 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8065 0.576 2.001 0.6325 ;
              RECT  1.923 0.417 2.001 0.6325 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.919 0.636 0.9615 0.951 ;
              RECT  0.919 0.3745 0.9615 0.4595 ;
              RECT  0.887 0.417 0.9295 0.6785 ;
              RECT  0.629 0.523 0.9295 0.5655 ;
              RECT  0.629 0.3815 0.6715 0.951 ;
              RECT  0.042 0.4735 0.6715 0.516 ;
              RECT  0.339 0.3815 0.3815 0.951 ;
              RECT  0.042 0.424 0.0985 0.516 ;
              RECT  0.049 0.3815 0.0985 0.516 ;
              RECT  0.049 0.3815 0.0915 0.951 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END SDFFHQX8

MACRO MDFFHQX2
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.212 0.3815 0.2545 0.9435 ;
              RECT  0.1835 0.5585 0.2545 0.6505 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.56 0.576 3.652 0.6325 ;
              RECT  3.5955 0.3535 3.638 0.6325 ;
              RECT  2.966 0.3535 3.638 0.3955 ;
              RECT  3.553 0.576 3.652 0.6185 ;
              RECT  3.1395 0.3535 3.224 0.4735 ;
              RECT  2.966 0.3535 3.0085 0.622 ;
        END
    END S0
    PIN D1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.295 0.555 3.4825 0.689 ;
              RECT  3.4255 0.4665 3.4825 0.689 ;
        END
    END D1
    PIN D0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7255 0.456 2.782 0.569 ;
              RECT  2.588 0.456 2.782 0.516 ;
              RECT  2.588 0.3535 2.6445 0.516 ;
        END
    END D0
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6645 0.576 0.721 ;
              RECT  0.449 0.629 0.576 0.721 ;
              RECT  0.325 0.6645 0.3815 0.788 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END MDFFHQX2

MACRO MX3X4
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.654 0.721 0.6965 0.997 ;
              RECT  0.654 0.2685 0.6965 0.3535 ;
              RECT  0.325 0.424 0.6645 0.4665 ;
              RECT  0.364 0.721 0.6965 0.7635 ;
              RECT  0.622 0.311 0.6645 0.4665 ;
              RECT  0.364 0.3675 0.4065 0.997 ;
              RECT  0.325 0.424 0.4065 0.516 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.107 0.728 2.503 0.7845 ;
              RECT  2.4465 0.6925 2.503 0.7845 ;
              RECT  2.107 0.7 2.1635 0.7845 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.2765 0.4735 2.503 0.53 ;
              RECT  2.305 0.4735 2.3615 0.6575 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.739 0.3425 1.796 0.6965 ;
        END
    END B
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.3425 1.6545 0.6965 ;
        END
    END S1
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.537 0.997 0.5935 ;
              RECT  0.8905 0.537 0.9475 0.841 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END MX3X4

MACRO MX2X2
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.424 1.23 0.516 ;
              RECT  1.0605 0.424 1.23 0.4665 ;
              RECT  1.0605 0.3005 1.103 0.781 ;
              RECT  1.0355 0.7385 1.078 1.0145 ;
              RECT  1.0355 0.258 1.078 0.3425 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8625 0.576 0.9895 0.6325 ;
              RECT  0.8625 0.576 0.919 0.859 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.311 0.675 0.438 0.7315 ;
              RECT  0.325 0.449 0.3815 0.7315 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.8025 0.5655 0.859 ;
              RECT  0.509 0.6575 0.5655 0.859 ;
              RECT  0.1835 0.6925 0.24 0.859 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END MX2X2

MACRO NAND4BBX4
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7255 0.3535 3.058 0.3955 ;
              RECT  3.0155 0.2965 3.058 0.3955 ;
              RECT  2.9235 0.767 2.966 0.965 ;
              RECT  0.894 0.767 2.966 0.8095 ;
              RECT  2.7255 0.2965 2.768 0.8095 ;
              RECT  2.6335 0.767 2.676 0.965 ;
              RECT  2.344 0.767 2.386 0.965 ;
              RECT  2.054 0.767 2.0965 0.965 ;
              RECT  1.764 0.767 1.8065 0.965 ;
              RECT  1.474 0.767 1.5165 0.965 ;
              RECT  1.184 0.767 1.2265 0.965 ;
              RECT  0.894 0.7105 1.1065 0.8095 ;
              RECT  0.894 0.7105 0.9365 0.965 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.5985 0.4595 2.655 0.6965 ;
              RECT  2.588 0.3535 2.6445 0.516 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.008 0.523 2.22 0.6965 ;
              RECT  2.008 0.4985 2.0645 0.6965 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.537 0.3815 0.8905 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.537 0.24 0.8905 ;
        END
    END BN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END NAND4BBX4

MACRO BMXIX2
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN PPN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8705 0.3815 2.927 0.912 ;
        END
    END PPN
    PIN X2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.588 0.371 2.6445 0.7245 ;
        END
    END X2
    PIN M1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2585 0.576 1.612 0.6325 ;
        END
    END M1
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.873 0.463 1.018 0.6325 ;
              RECT  0.8235 0.622 0.9295 0.6785 ;
        END
    END A
    PIN S
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.403 0.9755 1.4175 1.018 ;
              RECT  0.403 0.7315 0.445 1.018 ;
              RECT  0.357 0.7315 0.445 0.774 ;
              RECT  0.3075 0.7105 0.3995 0.767 ;
              RECT  0.3145 0.7035 0.3995 0.767 ;
        END
    END S
    PIN M0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.47 0.576 0.5265 0.661 ;
              RECT  0.166 0.576 0.5265 0.6325 ;
              RECT  0.1765 0.576 0.233 0.661 ;
        END
    END M0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END BMXIX2

MACRO AOI2BB1X2
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.318 0.636 0.3605 ;
              RECT  0.5935 0.2615 0.636 0.3605 ;
              RECT  0.449 0.7385 0.491 1.011 ;
              RECT  0.0565 0.7385 0.491 0.781 ;
              RECT  0.304 0.2615 0.346 0.3605 ;
              RECT  0.0565 0.318 0.0985 0.781 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2545 0.4985 0.6785 0.555 ;
              RECT  0.325 0.4985 0.3815 0.6505 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7915 0.424 0.8485 0.629 ;
              RECT  0.7495 0.318 0.806 0.516 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.3995 1.0885 0.753 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END AOI2BB1X2

MACRO TBUFX6
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.623 0.3745 2.9555 0.417 ;
              RECT  2.913 0.318 2.9555 0.417 ;
              RECT  2.8775 0.3745 2.92 0.912 ;
              RECT  2.4465 0.636 2.92 0.6785 ;
              RECT  2.623 0.318 2.6655 0.417 ;
              RECT  2.588 0.636 2.63 0.912 ;
              RECT  2.4465 0.5585 2.503 0.6785 ;
              RECT  2.298 0.7 2.489 0.742 ;
              RECT  2.4465 0.41 2.489 0.742 ;
              RECT  2.333 0.41 2.489 0.4525 ;
              RECT  2.333 0.318 2.3755 0.4525 ;
              RECT  2.298 0.7 2.3405 0.912 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.001 0.187 2.1425 0.2295 ;
              RECT  0.94 0.1905 2.0435 0.233 ;
              RECT  0.417 0.608 0.9825 0.6505 ;
              RECT  0.94 0.1905 0.9825 0.6505 ;
              RECT  0.449 0.576 0.5405 0.6505 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.827 0.4525 0.8695 0.537 ;
              RECT  0.1835 0.463 0.8695 0.5055 ;
              RECT  0.6115 0.463 0.6965 0.5335 ;
              RECT  0.1555 0.608 0.24 0.6505 ;
              RECT  0.1835 0.463 0.24 0.6505 ;
        END
    END OE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END TBUFX6

MACRO TBUFX12
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.43 0.608 4.472 0.993 ;
              RECT  3.012 0.608 4.472 0.6505 ;
              RECT  3.7685 0.35 4.391 0.392 ;
              RECT  4.3485 0.293 4.391 0.392 ;
              RECT  4.14 0.35 4.1825 0.993 ;
              RECT  4.0585 0.293 4.101 0.392 ;
              RECT  3.85 0.608 3.8925 0.993 ;
              RECT  3.7685 0.293 3.811 0.392 ;
              RECT  3.56 0.608 3.6025 0.993 ;
              RECT  3.189 0.35 3.521 0.392 ;
              RECT  3.4785 0.293 3.521 0.392 ;
              RECT  3.27 0.35 3.3125 0.993 ;
              RECT  3.189 0.293 3.231 0.392 ;
              RECT  3.012 0.5585 3.0685 0.6505 ;
              RECT  3.012 0.35 3.0545 0.7635 ;
              RECT  2.98 0.721 3.0225 0.993 ;
              RECT  2.899 0.35 3.0545 0.392 ;
              RECT  2.899 0.293 2.9415 0.392 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.6685 0.569 2.6725 0.6115 ;
              RECT  2.63 0.5265 2.6725 0.6115 ;
              RECT  1.6685 0.456 1.711 0.6115 ;
              RECT  1.46 0.456 1.711 0.4985 ;
              RECT  1.46 0.205 1.5025 0.4985 ;
              RECT  1.1735 0.205 1.5025 0.247 ;
              RECT  0.905 0.4345 1.216 0.477 ;
              RECT  1.1735 0.205 1.216 0.477 ;
              RECT  0.905 0.2085 0.9475 0.477 ;
              RECT  0.636 0.2085 0.9475 0.251 ;
              RECT  0.3815 0.569 0.6785 0.6115 ;
              RECT  0.636 0.2085 0.6785 0.6115 ;
              RECT  0.449 0.569 0.5405 0.6325 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2545 0.4415 0.5655 0.4985 ;
              RECT  0.509 0.4135 0.5655 0.4985 ;
              RECT  0.2545 0.4415 0.311 0.5515 ;
        END
    END OE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END TBUFX12

MACRO NAND3X1
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.8485 0.6645 1.0535 ;
              RECT  0.608 0.311 0.6505 1.0535 ;
              RECT  0.3005 0.8485 0.6645 0.8905 ;
              RECT  0.5265 0.311 0.6505 0.3535 ;
              RECT  0.5265 0.2685 0.569 0.3535 ;
              RECT  0.3005 0.8485 0.3425 1.0465 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.424 0.523 0.7775 ;
        END
    END C
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.339 0.3955 0.629 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END NAND3X1

MACRO DFFSRHQX2
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.293 0.8445 0.3995 0.9015 ;
              RECT  0.293 0.3815 0.3355 0.919 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.426 0.424 4.483 0.7775 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.9845 0.4415 4.076 0.4985 ;
              RECT  3.825 0.544 4.041 0.601 ;
              RECT  3.9845 0.4415 4.041 0.601 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.775 0.9825 3.058 1.025 ;
              RECT  2.775 0.8485 2.8175 1.025 ;
              RECT  2.5065 0.8485 2.8175 0.8905 ;
              RECT  1.7885 0.905 2.549 0.9475 ;
              RECT  2.5065 0.8485 2.549 0.9475 ;
              RECT  1.7885 0.8485 1.831 0.9475 ;
              RECT  1.4315 0.8485 1.831 0.8905 ;
              RECT  1.2055 0.8625 1.474 0.905 ;
              RECT  1.2055 0.7105 1.248 0.905 ;
              RECT  1.202 0.5865 1.2445 0.767 ;
              RECT  1.156 0.7105 1.248 0.767 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.5865 1.085 0.643 ;
              RECT  0.8905 0.5865 0.9475 0.8025 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END DFFSRHQX2

MACRO NAND4BBX1
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9085 0.2155 0.951 0.767 ;
              RECT  0.905 0.6925 0.9475 1.0465 ;
              RECT  0.4345 0.2155 0.951 0.258 ;
              RECT  0.601 0.8485 0.9475 0.8905 ;
              RECT  0.8905 0.6925 0.9475 0.8905 ;
              RECT  0.601 0.8485 0.643 1.0465 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3425 0.4415 0.5195 0.4985 ;
              RECT  0.3075 0.576 0.3995 0.6395 ;
              RECT  0.3425 0.4415 0.3995 0.6395 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.59 0.5585 0.6645 0.7775 ;
              RECT  0.59 0.4415 0.647 0.7775 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.191 0.548 1.248 0.866 ;
              RECT  1.156 0.576 1.248 0.6325 ;
              RECT  1.184 0.548 1.248 0.6325 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.622 0.1235 0.7315 ;
              RECT  0.042 0.424 0.0985 0.7315 ;
              RECT  0.021 0.424 0.0985 0.516 ;
        END
    END BN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END NAND4BBX1

MACRO DFFHQX1
    CLASS CORE ;
    SIZE 2.5455 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.081 0.3675 0.1235 1.0465 ;
              RECT  0.042 0.424 0.1235 0.516 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.199 0.5195 2.3825 0.7455 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.537 0.3815 0.8905 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.5455 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.5455 0.042 ;
        END
    END VSS
END DFFHQX1

MACRO SEDFFTRXL
    CLASS CORE ;
    SIZE 5.6565 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.8005 0.5265 3.917 0.583 ;
              RECT  3.8605 0.2755 3.917 0.583 ;
              RECT  3.8005 0.5265 3.857 0.735 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.2895 0.1165 0.449 ;
              RECT  0.042 0.2895 0.0985 0.721 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.4305 0.5195 5.487 0.7495 ;
              RECT  5.416 0.6925 5.473 0.859 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.907 0.544 5.229 0.601 ;
              RECT  4.974 0.544 5.066 0.6325 ;
        END
    END E
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1045 0.661 4.292 0.7175 ;
              RECT  4.1435 0.661 4.2 0.8835 ;
        END
    END RN
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.952 0.5265 3.0935 0.668 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.3195 0.4135 3.362 0.4985 ;
              RECT  2.839 0.4135 3.362 0.456 ;
              RECT  2.7115 0.4415 2.881 0.4985 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.2765 0.523 2.4145 0.6325 ;
              RECT  2.2765 0.5195 2.333 0.7915 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.6565 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.6565 0.042 ;
        END
    END VSS
END SEDFFTRXL

MACRO TLATNTSCAX6
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.309 0.537 3.3515 0.9685 ;
              RECT  3.309 0.247 3.3515 0.4665 ;
              RECT  3.277 0.424 3.3195 0.5795 ;
              RECT  2.729 0.537 3.3515 0.5795 ;
              RECT  3.019 0.247 3.0615 0.9685 ;
              RECT  2.729 0.537 2.786 0.6505 ;
              RECT  2.729 0.247 2.7715 0.9685 ;
        END
    END ECK
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.318 0.523 0.6715 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.318 0.3815 0.6715 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0245 0.576 0.141 0.6325 ;
              RECT  0.0565 0.339 0.141 0.6325 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END TLATNTSCAX6

MACRO SDFFRHQX4
    CLASS CORE ;
    SIZE 5.091 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.833 0.4415 4.9245 0.4985 ;
              RECT  4.833 0.35 4.8755 0.4985 ;
              RECT  4.3695 0.35 4.8755 0.392 ;
              RECT  4.3695 0.35 4.4545 0.47 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.5675 0.5585 4.762 0.6785 ;
              RECT  4.7055 0.463 4.762 0.6785 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1115 0.4415 4.168 0.622 ;
              RECT  3.9385 0.4415 4.168 0.4985 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.503 0.5975 2.7785 0.6395 ;
              RECT  2.7365 0.537 2.7785 0.6395 ;
              RECT  2.503 0.2365 2.5455 0.6395 ;
              RECT  1.2125 0.2365 2.5455 0.279 ;
              RECT  1.559 0.2365 1.6015 0.5265 ;
              RECT  1.1735 0.424 1.255 0.5335 ;
              RECT  1.2125 0.2365 1.255 0.5335 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.484 0.24 0.8375 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.866 0.3885 0.9615 0.431 ;
              RECT  0.8235 0.6785 0.9085 0.721 ;
              RECT  0.866 0.3885 0.9085 0.721 ;
              RECT  0.608 0.424 0.9085 0.4665 ;
              RECT  0.491 0.6785 0.6645 0.721 ;
              RECT  0.622 0.3675 0.6645 0.721 ;
              RECT  0.608 0.3675 0.6645 0.516 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.091 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.091 0.042 ;
        END
    END VSS
END SDFFRHQX4

MACRO NAND2XL
    CLASS CORE ;
    SIZE 0.5655 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.212 0.806 0.4945 0.8485 ;
              RECT  0.4525 0.339 0.4945 0.8485 ;
              RECT  0.325 0.339 0.4945 0.3815 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.1835 0.6505 ;
              RECT  0.127 0.4525 0.1835 0.6505 ;
              RECT  0.042 0.5585 0.0985 0.721 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2545 0.5585 0.3815 0.735 ;
              RECT  0.279 0.4525 0.3815 0.735 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.5655 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.5655 0.042 ;
        END
    END VSS
END NAND2XL

MACRO TBUFX4
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7355 0.6645 1.778 0.94 ;
              RECT  1.4565 0.6645 1.778 0.707 ;
              RECT  1.375 0.346 1.7075 0.3885 ;
              RECT  1.665 0.2895 1.7075 0.3885 ;
              RECT  1.4565 0.5585 1.513 0.707 ;
              RECT  1.4565 0.346 1.499 0.813 ;
              RECT  1.446 0.7705 1.488 0.94 ;
              RECT  1.375 0.2895 1.4175 0.3885 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0745 0.431 1.1595 0.4735 ;
              RECT  1.117 0.1975 1.1595 0.4735 ;
              RECT  0.59 0.1975 1.1595 0.24 ;
              RECT  0.59 0.4415 0.682 0.4985 ;
              RECT  0.3145 0.5865 0.6325 0.629 ;
              RECT  0.59 0.1975 0.6325 0.629 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.187 0.4595 0.5195 0.516 ;
              RECT  0.325 0.424 0.3815 0.516 ;
              RECT  0.187 0.4595 0.2435 0.544 ;
        END
    END OE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END TBUFX4

MACRO AOI2BB2XL
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.322 0.576 1.534 0.6325 ;
              RECT  1.322 0.463 1.3785 0.661 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0815 0.4415 1.138 0.59 ;
              RECT  0.8765 0.4415 1.138 0.4985 ;
        END
    END B1
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3355 0.325 0.3995 0.643 ;
              RECT  0.3075 0.325 0.3995 0.3815 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.4525 0.24 0.806 ;
        END
    END A1N
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.209 0.7315 1.294 0.774 ;
              RECT  1.209 0.3285 1.2515 0.774 ;
              RECT  0.7635 0.3285 1.2515 0.371 ;
              RECT  0.7495 0.424 0.806 0.516 ;
              RECT  0.7635 0.3285 0.806 0.516 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END AOI2BB2XL

MACRO SDFFNSRXL
    CLASS CORE ;
    SIZE 5.6565 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.834 0.8305 0.919 ;
              RECT  0.774 0.2615 0.8305 0.346 ;
              RECT  0.608 0.827 0.788 0.919 ;
              RECT  0.7315 0.2895 0.788 0.919 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.721 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.3985 0.4415 5.4905 0.4985 ;
              RECT  5.4055 0.4415 5.448 0.5265 ;
              RECT  5.0095 0.47 5.448 0.5125 ;
              RECT  5.0095 0.47 5.1685 0.555 ;
              RECT  5.0095 0.47 5.052 0.742 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.3985 0.6045 5.4905 0.767 ;
              RECT  5.243 0.6045 5.4905 0.661 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.6065 0.7105 4.826 0.767 ;
              RECT  4.6915 0.576 4.7835 0.767 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.3945 0.7105 4.536 0.767 ;
              RECT  4.3945 0.583 4.536 0.6395 ;
              RECT  4.3945 0.583 4.451 0.767 ;
        END
    END CKN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.0755 0.9225 3.3975 0.965 ;
              RECT  3.0755 0.8305 3.118 0.965 ;
              RECT  1.612 0.8305 3.118 0.873 ;
              RECT  1.612 0.6925 1.6545 0.873 ;
              RECT  1.598 0.583 1.64 0.7845 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0145 0.53 1.1065 0.7915 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.6565 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.6565 0.042 ;
        END
    END VSS
END SDFFNSRXL

MACRO ADDFHX1
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN CI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5625 0.3885 2.39 0.431 ;
              RECT  1.1345 0.346 1.605 0.3885 ;
              RECT  1.1345 0.3075 1.248 0.3885 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.588 0.502 2.6725 0.5585 ;
              RECT  2.588 0.502 2.6445 0.6505 ;
              RECT  1.354 0.502 2.6725 0.544 ;
              RECT  0.622 0.463 1.3965 0.5055 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4745 0.615 2.517 0.7 ;
              RECT  1.2405 0.615 2.517 0.6575 ;
              RECT  0.8025 0.576 1.283 0.6185 ;
              RECT  1.156 0.615 2.517 0.6325 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2435 0.6505 0.286 0.912 ;
              RECT  0.042 0.424 0.286 0.4665 ;
              RECT  0.2435 0.3675 0.286 0.4665 ;
              RECT  0.0565 0.6505 0.286 0.6925 ;
              RECT  0.0565 0.424 0.0985 0.6925 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.899 0.424 3.0685 0.516 ;
              RECT  2.899 0.3815 2.9415 0.912 ;
        END
    END S
END ADDFHX1

MACRO SDFFRHQX1
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.067 0.318 0.1235 0.997 ;
              RECT  0.042 0.424 0.1235 0.516 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.783 0.456 3.825 0.5405 ;
              RECT  3.7015 0.4415 3.7935 0.4985 ;
              RECT  3.2385 0.456 3.825 0.4985 ;
              RECT  3.2385 0.456 3.2805 0.707 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4715 0.569 3.712 0.6255 ;
              RECT  3.4715 0.569 3.652 0.7385 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.998 0.424 3.0545 0.615 ;
              RECT  2.8705 0.424 3.0545 0.4805 ;
              RECT  2.8705 0.424 2.927 0.516 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0145 0.576 1.163 0.7245 ;
              RECT  0.933 0.544 1.071 0.601 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.4875 0.3815 0.841 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END SDFFRHQX1

MACRO CLKMX2X3
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.534 0.608 1.5765 0.965 ;
              RECT  1.276 0.3675 1.5765 0.41 ;
              RECT  1.534 0.311 1.5765 0.41 ;
              RECT  1.276 0.608 1.5765 0.6505 ;
              RECT  1.276 0.5585 1.3715 0.6505 ;
              RECT  1.276 0.332 1.3185 0.7455 ;
              RECT  1.2445 0.7035 1.2865 0.965 ;
              RECT  1.223 0.332 1.3185 0.3745 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0145 0.576 1.2055 0.6325 ;
              RECT  1.0145 0.5585 1.071 0.7775 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.449 0.5585 0.562 0.7175 ;
              RECT  0.311 0.5585 0.562 0.615 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6325 0.5935 0.7175 0.636 ;
              RECT  0.1975 0.788 0.675 0.8305 ;
              RECT  0.6325 0.5935 0.675 0.8305 ;
              RECT  0.1975 0.5585 0.24 0.8305 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END CLKMX2X3

MACRO EDFFTRX1
    CLASS CORE ;
    SIZE 5.091 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6715 0.357 0.714 0.4525 ;
              RECT  0.6645 0.424 0.707 0.82 ;
              RECT  0.608 0.424 0.707 0.516 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.912 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.762 0.6925 4.907 0.7845 ;
              RECT  4.8505 0.5195 4.907 0.7845 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4085 0.5585 4.5005 0.6325 ;
              RECT  4.122 0.5585 4.5005 0.615 ;
        END
    END E
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4365 0.5585 3.493 0.806 ;
              RECT  3.33 0.5585 3.493 0.615 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.898 0.4945 0.9545 0.7495 ;
              RECT  0.8905 0.6925 0.9475 0.841 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.091 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.091 0.042 ;
        END
    END VSS
END EDFFTRX1

MACRO DFFX1
    CLASS CORE ;
    SIZE 2.9695 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.622 0.3815 0.6645 0.9475 ;
              RECT  0.608 0.3815 0.6645 0.516 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1445 0.3815 0.2015 0.912 ;
              RECT  0.042 0.424 0.2015 0.516 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.471 0.7105 2.7435 0.767 ;
              RECT  2.57 0.629 2.6265 0.767 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.852 0.5515 0.9085 0.636 ;
              RECT  0.7495 0.6925 0.905 0.8025 ;
              RECT  0.8485 0.5795 0.905 0.8025 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.9695 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.9695 0.042 ;
        END
    END VSS
END DFFX1

MACRO MDFFHQX8
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.483 0.4415 4.525 0.5265 ;
              RECT  4.4085 0.4415 4.525 0.4985 ;
              RECT  3.977 0.456 4.525 0.4985 ;
              RECT  3.9135 0.491 4.0195 0.5335 ;
              RECT  3.9135 0.491 3.956 0.682 ;
        END
    END S0
    PIN D1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.147 0.569 4.412 0.6255 ;
              RECT  4.147 0.569 4.359 0.714 ;
        END
    END D1
    PIN D0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.673 0.5585 3.7295 0.7175 ;
              RECT  3.5775 0.5585 3.7295 0.6505 ;
              RECT  3.5775 0.4595 3.6345 0.6505 ;
        END
    END D0
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8065 0.576 2.001 0.6325 ;
              RECT  1.923 0.417 2.001 0.6325 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.919 0.636 0.9615 0.951 ;
              RECT  0.919 0.3745 0.9615 0.4595 ;
              RECT  0.887 0.417 0.9295 0.6785 ;
              RECT  0.629 0.523 0.9295 0.5655 ;
              RECT  0.629 0.3815 0.6715 0.951 ;
              RECT  0.042 0.4735 0.6715 0.516 ;
              RECT  0.339 0.3815 0.3815 0.951 ;
              RECT  0.042 0.424 0.0985 0.516 ;
              RECT  0.049 0.3815 0.0985 0.516 ;
              RECT  0.049 0.3815 0.0915 0.951 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END MDFFHQX8

MACRO CLKAND2X8
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.2485 0.668 2.291 0.9825 ;
              RECT  2.1775 0.3605 2.273 0.403 ;
              RECT  1.3785 0.668 2.291 0.7105 ;
              RECT  2.1635 0.5585 2.22 0.7105 ;
              RECT  1.361 0.371 2.2095 0.4135 ;
              RECT  2.1635 0.371 2.206 0.7105 ;
              RECT  1.9585 0.668 2.001 0.9825 ;
              RECT  1.8985 0.3605 1.983 0.4135 ;
              RECT  1.6685 0.668 1.711 0.9825 ;
              RECT  1.6085 0.3605 1.6935 0.4135 ;
              RECT  1.3785 0.668 1.421 0.9825 ;
              RECT  1.3185 0.3605 1.4035 0.403 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.431 0.576 0.965 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.092 0.463 1.1345 0.548 ;
              RECT  0.166 0.463 1.1345 0.5055 ;
              RECT  0.166 0.4415 0.258 0.5055 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END CLKAND2X8

MACRO CLKINVX20
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.5735 0.6395 2.616 0.9615 ;
              RECT  0.774 0.6505 2.616 0.6925 ;
              RECT  0.194 0.424 2.556 0.4665 ;
              RECT  2.5135 0.251 2.556 0.4665 ;
              RECT  2.4465 0.5585 2.503 0.6925 ;
              RECT  2.333 0.424 2.3755 0.6925 ;
              RECT  2.2235 0.6505 2.266 0.9615 ;
              RECT  2.2235 0.251 2.266 0.4665 ;
              RECT  1.9335 0.6505 1.976 0.9615 ;
              RECT  1.9335 0.251 1.976 0.4665 ;
              RECT  1.644 0.6505 1.686 0.9615 ;
              RECT  1.644 0.251 1.686 0.4665 ;
              RECT  1.354 0.6505 1.3965 0.9615 ;
              RECT  1.354 0.251 1.3965 0.4665 ;
              RECT  1.064 0.6505 1.1065 0.9615 ;
              RECT  1.064 0.251 1.1065 0.4665 ;
              RECT  0.774 0.6505 0.8165 0.9615 ;
              RECT  0.774 0.251 0.8165 0.4665 ;
              RECT  0.194 0.7635 0.8165 0.806 ;
              RECT  0.484 0.6505 0.5265 0.9615 ;
              RECT  0.484 0.251 0.5265 0.4665 ;
              RECT  0.194 0.6505 0.2365 0.9615 ;
              RECT  0.194 0.251 0.2365 0.4665 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.226 0.537 2.1955 0.5795 ;
              RECT  0.3075 0.537 0.3995 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END CLKINVX20

MACRO OA21XL
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.403 0.9755 0.4595 ;
              RECT  0.742 0.4595 0.9475 0.516 ;
              RECT  0.742 0.4595 0.799 0.8375 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3955 0.24 0.7495 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.1555 0.523 0.509 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END OA21XL

MACRO OAI211X2
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.382 0.3215 1.506 0.364 ;
              RECT  0.905 0.449 1.4245 0.491 ;
              RECT  1.382 0.3215 1.4245 0.491 ;
              RECT  1.237 0.7495 1.2795 0.951 ;
              RECT  0.4525 0.7495 1.2795 0.7915 ;
              RECT  0.9475 0.7495 0.9895 0.951 ;
              RECT  0.8905 0.6925 0.9475 0.7915 ;
              RECT  0.905 0.449 0.9475 0.7915 ;
              RECT  0.4525 0.7495 0.4945 0.951 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.576 0.5265 0.6325 ;
              RECT  0.325 0.576 0.3815 0.7845 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.449 0.689 0.5055 ;
              RECT  0.1975 0.449 0.2545 0.622 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.018 0.562 1.3115 0.6785 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.5585 1.6545 0.6855 ;
              RECT  1.4955 0.5585 1.6545 0.6325 ;
              RECT  1.4955 0.4345 1.552 0.6325 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END OAI211X2

MACRO TBUFX2
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.2615 1.3715 0.905 ;
              RECT  1.2975 0.2615 1.3715 0.346 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9895 0.4875 1.0745 0.53 ;
              RECT  0.4985 0.806 1.032 0.8485 ;
              RECT  0.9895 0.4875 1.032 0.8485 ;
              RECT  0.4985 0.576 0.5405 0.8485 ;
              RECT  0.449 0.576 0.5405 0.6325 ;
              RECT  0.392 0.569 0.491 0.6115 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.4415 0.5405 0.4985 ;
              RECT  0.205 0.4415 0.286 0.5265 ;
        END
    END OE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END TBUFX2

MACRO DFFSRX4
    CLASS CORE ;
    SIZE 5.798 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.9175 0.318 5.335 0.3605 ;
              RECT  5.25 0.647 5.2925 0.9225 ;
              RECT  4.939 0.647 5.2925 0.689 ;
              RECT  4.992 0.318 5.0485 0.689 ;
              RECT  4.939 0.647 4.9815 0.9225 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.253 0.311 4.67 0.3535 ;
              RECT  4.5925 0.647 4.635 0.9225 ;
              RECT  4.285 0.647 4.635 0.689 ;
              RECT  4.299 0.311 4.3415 0.689 ;
              RECT  4.285 0.424 4.327 0.9225 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.259 0.576 2.4815 0.6325 ;
              RECT  2.287 0.445 2.4815 0.6325 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.9655 0.576 2.188 0.6325 ;
              RECT  2.0045 0.445 2.188 0.6325 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3145 0.7105 0.5405 0.767 ;
              RECT  0.41 0.583 0.5405 0.767 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.445 0.24 0.799 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.798 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.798 0.042 ;
        END
    END VSS
END DFFSRX4

MACRO ADDHX1
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.022 0.3885 2.0785 0.6855 ;
              RECT  1.9865 0.629 2.0435 0.912 ;
              RECT  1.9865 0.3605 2.0435 0.445 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1235 0.293 0.166 1.039 ;
              RECT  0.042 0.424 0.166 0.516 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.4415 0.742 0.5795 ;
              RECT  0.47 0.4415 0.742 0.4985 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.039 0.265 1.3505 0.3075 ;
              RECT  1.039 0.2015 1.0815 0.3075 ;
              RECT  0.424 0.2015 1.0815 0.2435 ;
              RECT  0.3145 0.3285 0.4665 0.371 ;
              RECT  0.424 0.2015 0.4665 0.371 ;
              RECT  0.3075 0.4415 0.3995 0.4985 ;
              RECT  0.3145 0.3285 0.3995 0.4985 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END ADDHX1

MACRO EDFFXL
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.8605 0.5585 3.917 0.8095 ;
              RECT  3.8675 0.293 3.917 0.8095 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.403 3.21 0.5655 ;
              RECT  3.1465 0.53 3.203 0.721 ;
              RECT  3.125 0.403 3.21 0.4595 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8705 0.5585 2.927 0.6505 ;
              RECT  2.4285 0.8905 2.899 0.933 ;
              RECT  2.8565 0.608 2.899 0.933 ;
              RECT  2.2415 0.993 2.471 1.0355 ;
              RECT  2.4285 0.4985 2.471 1.0355 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.662 0.5335 2.786 0.82 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5405 0.24 0.894 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END EDFFXL

MACRO OAI21XL
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4525 0.8485 0.6645 0.8905 ;
              RECT  0.608 0.6925 0.6645 0.8905 ;
              RECT  0.608 0.311 0.6505 0.8905 ;
              RECT  0.5335 0.311 0.6505 0.3535 ;
              RECT  0.5335 0.2685 0.576 0.3535 ;
              RECT  0.4525 0.8485 0.4945 0.979 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.537 0.0985 0.8905 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5655 0.3815 0.919 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.424 0.523 0.7775 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END OAI21XL

MACRO MX2X8
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3085 0.35 2.351 1.0145 ;
              RECT  1.4385 0.7 2.351 0.742 ;
              RECT  1.7605 0.392 2.351 0.4345 ;
              RECT  1.9975 0.3815 2.082 0.4345 ;
              RECT  2.0185 0.7 2.061 1.0145 ;
              RECT  1.7075 0.3815 1.7925 0.424 ;
              RECT  1.7285 0.7 1.771 1.0145 ;
              RECT  1.4565 0.6925 1.513 0.7845 ;
              RECT  1.4565 0.3745 1.499 0.7845 ;
              RECT  1.4385 0.7 1.481 1.0145 ;
              RECT  1.414 0.3745 1.499 0.417 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.601 1.23 0.841 ;
              RECT  1.0605 0.601 1.23 0.6575 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.449 0.5055 0.5655 0.767 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.636 0.6115 0.721 0.654 ;
              RECT  0.3355 0.8375 0.6785 0.88 ;
              RECT  0.636 0.6115 0.6785 0.88 ;
              RECT  0.3355 0.675 0.378 0.88 ;
              RECT  0.1835 0.675 0.378 0.7845 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END MX2X8

MACRO CLKMX2X6
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7355 0.654 1.778 0.986 ;
              RECT  1.718 0.166 1.7605 0.385 ;
              RECT  1.704 0.3425 1.7465 0.6965 ;
              RECT  1.17 0.424 1.7465 0.4665 ;
              RECT  1.446 0.424 1.488 0.986 ;
              RECT  1.428 0.166 1.4705 0.4665 ;
              RECT  1.17 0.424 1.23 0.622 ;
              RECT  1.17 0.251 1.2125 0.622 ;
              RECT  1.156 0.5865 1.1985 0.986 ;
              RECT  1.138 0.2085 1.1805 0.293 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.477 0.9475 0.8305 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.4665 0.7035 ;
              RECT  0.41 0.4345 0.4665 0.7035 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.774 0.5935 0.8305 ;
              RECT  0.537 0.647 0.5935 0.8305 ;
              RECT  0.1835 0.647 0.2545 0.7845 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END CLKMX2X6

MACRO EDFFTRX4
    CLASS CORE ;
    SIZE 5.9395 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.1475 0.6575 5.579 0.7 ;
              RECT  5.1475 0.364 5.4835 0.4065 ;
              RECT  5.441 0.3075 5.4835 0.4065 ;
              RECT  5.1475 0.3075 5.1935 0.4065 ;
              RECT  5.1475 0.3075 5.19 0.7 ;
              RECT  5.1335 0.5585 5.19 0.6505 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.497 0.6575 4.914 0.7 ;
              RECT  4.571 0.364 4.9035 0.4065 ;
              RECT  4.861 0.3075 4.9035 0.4065 ;
              RECT  4.709 0.5585 4.7655 0.7 ;
              RECT  4.709 0.364 4.7515 0.7 ;
              RECT  4.571 0.3075 4.6135 0.4065 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.825 0.622 4.002 0.6785 ;
              RECT  3.843 0.576 4.002 0.6785 ;
              RECT  3.843 0.445 3.9985 0.6785 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.895 0.576 2.199 0.6325 ;
              RECT  1.895 0.576 2.0965 0.682 ;
        END
    END RN
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9225 0.608 1.025 0.6505 ;
              RECT  0.449 0.859 0.965 0.9015 ;
              RECT  0.9225 0.608 0.965 0.9015 ;
              RECT  0.449 0.8445 0.5405 0.9015 ;
              RECT  0.4985 0.569 0.5405 0.9015 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5585 0.4275 0.6505 ;
              RECT  0.371 0.5195 0.4275 0.6505 ;
              RECT  0.1835 0.5585 0.24 0.6855 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.9395 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.9395 0.042 ;
        END
    END VSS
END EDFFTRX4

MACRO NOR2BX1
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.251 0.2615 0.293 0.346 ;
              RECT  0.0565 0.318 0.2615 0.3605 ;
              RECT  0.219 0.304 0.293 0.346 ;
              RECT  0.1765 0.8555 0.219 0.94 ;
              RECT  0.0565 0.8555 0.219 0.898 ;
              RECT  0.0565 0.318 0.0985 0.898 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.53 0.5405 0.7105 ;
              RECT  0.311 0.576 0.5405 0.6325 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.24 0.7845 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END NOR2BX1

MACRO SDFFSRX1
    CLASS CORE ;
    SIZE 5.2325 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6325 0.5865 0.675 1.011 ;
              RECT  0.6325 0.258 0.675 0.3425 ;
              RECT  0.622 0.311 0.6645 0.629 ;
              RECT  0.608 0.424 0.6645 0.516 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1695 0.3815 0.226 0.912 ;
              RECT  0.042 0.424 0.226 0.516 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.006 0.4415 5.0485 0.5265 ;
              RECT  4.4935 0.463 5.0485 0.5055 ;
              RECT  4.833 0.4415 5.0485 0.5055 ;
              RECT  4.7195 0.4205 4.762 0.5055 ;
              RECT  4.4935 0.463 4.536 0.707 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.6065 0.601 4.9355 0.6575 ;
              RECT  4.6915 0.576 4.9355 0.6575 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.956 0.576 4.3095 0.6325 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.0195 0.7035 4.3095 0.76 ;
              RECT  3.963 0.7105 4.076 0.767 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.747 0.9295 3.111 0.972 ;
              RECT  2.747 0.8165 2.7895 0.972 ;
              RECT  2.1105 0.8165 2.7895 0.859 ;
              RECT  2.1105 0.654 2.153 0.859 ;
              RECT  1.4385 0.654 2.153 0.6965 ;
              RECT  1.4385 0.576 1.5305 0.6965 ;
              RECT  1.4105 0.576 1.5305 0.6185 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.502 0.9475 0.8555 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.2325 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.2325 0.042 ;
        END
    END VSS
END SDFFSRX1

MACRO CLKAND2X2
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5655 0.424 0.6645 0.516 ;
              RECT  0.4985 0.5795 0.608 0.622 ;
              RECT  0.5655 0.2545 0.608 0.622 ;
              RECT  0.4985 0.2545 0.608 0.2965 ;
              RECT  0.4985 0.5795 0.5405 0.9475 ;
              RECT  0.4985 0.212 0.5405 0.2965 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.3815 0.7915 ;
              RECT  0.2825 0.4805 0.3425 0.7495 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.0985 0.912 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END CLKAND2X2

MACRO OAI22X1
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.59 0.41 0.682 0.4525 ;
              RECT  0.6395 0.3675 0.682 0.4525 ;
              RECT  0.59 0.41 0.6325 0.5725 ;
              RECT  0.4805 0.53 0.6325 0.5725 ;
              RECT  0.4805 0.53 0.523 1.032 ;
              RECT  0.4665 0.5585 0.523 0.6505 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.636 0.3955 0.8695 ;
              RECT  0.339 0.53 0.3955 0.8695 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.53 0.24 0.7845 ;
              RECT  0.0845 0.53 0.24 0.5865 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.523 0.806 0.8765 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.827 0.6645 0.9825 ;
              RECT  0.5935 0.643 0.6505 0.8695 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END OAI22X1

MACRO DFFSRX2
    CLASS CORE ;
    SIZE 5.6565 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.1335 0.403 5.271 0.4595 ;
              RECT  5.151 0.647 5.2075 0.9225 ;
              RECT  5.1335 0.403 5.19 0.7845 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.8645 0.3815 4.921 0.9225 ;
              RECT  4.8505 0.6925 4.921 0.7845 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.5395 0.7105 4.681 0.767 ;
              RECT  4.624 0.4985 4.681 0.767 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2975 0.576 1.4105 0.753 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.463 0.6715 0.721 0.728 ;
              RECT  0.463 0.576 0.682 0.728 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1095 0.325 0.166 0.576 ;
              RECT  0.042 0.325 0.166 0.3815 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.6565 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.6565 0.042 ;
        END
    END VSS
END DFFSRX2

MACRO OAI32X1
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.622 0.4595 0.8905 0.502 ;
              RECT  0.8485 0.311 0.8905 0.502 ;
              RECT  0.622 0.4595 0.6645 0.9615 ;
              RECT  0.608 0.5585 0.6645 0.6505 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3675 0.24 0.721 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5655 0.3815 0.919 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.5725 0.806 0.926 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4805 0.4595 0.537 0.735 ;
              RECT  0.4665 0.6925 0.523 0.799 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9615 0.3675 1.0885 0.516 ;
              RECT  0.9615 0.3675 1.018 0.6505 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END OAI32X1

MACRO TLATNCAX6
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8845 0.247 2.927 0.9755 ;
              RECT  2.305 0.53 2.927 0.5725 ;
              RECT  2.595 0.247 2.6375 0.9755 ;
              RECT  2.305 0.424 2.3615 0.5725 ;
              RECT  2.305 0.247 2.3475 0.9755 ;
        END
    END ECK
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.7105 0.5405 0.9435 ;
              RECT  0.424 0.7105 0.5405 0.767 ;
              RECT  0.424 0.6505 0.4805 0.767 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2965 0.5125 0.3535 0.735 ;
              RECT  0.166 0.548 0.3535 0.6325 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END TLATNCAX6

MACRO OA22XL
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1275 0.3005 1.17 1.004 ;
              RECT  1.032 0.9615 1.17 1.004 ;
              RECT  0.919 0.9825 1.0885 1.0535 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.537 0.806 0.8905 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.424 0.3955 0.7635 ;
              RECT  0.325 0.424 0.3955 0.516 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.509 0.4735 0.5655 0.7495 ;
              RECT  0.4665 0.6925 0.523 0.7845 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OA22XL

MACRO AND2X8
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.6685 0.6925 1.711 1.0075 ;
              RECT  1.598 0.339 1.6935 0.3815 ;
              RECT  0.799 0.6925 1.711 0.735 ;
              RECT  0.781 0.35 1.6295 0.392 ;
              RECT  1.4565 0.35 1.513 0.516 ;
              RECT  1.4565 0.35 1.499 0.735 ;
              RECT  1.3785 0.6925 1.421 1.0075 ;
              RECT  1.3185 0.339 1.4035 0.392 ;
              RECT  1.0885 0.6925 1.131 1.0075 ;
              RECT  1.0285 0.339 1.1135 0.392 ;
              RECT  0.799 0.6925 0.841 1.0075 ;
              RECT  0.7385 0.339 0.8235 0.3815 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.569 0.4275 0.7385 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4985 0.4415 0.555 0.5265 ;
              RECT  0.0245 0.4415 0.555 0.4985 ;
              RECT  0.152 0.4415 0.2365 0.502 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END AND2X8

MACRO TLATNX4
    CLASS CORE ;
    SIZE 3.6765 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8735 0.364 2.2485 0.4065 ;
              RECT  2.206 0.3215 2.2485 0.4065 ;
              RECT  2.0785 0.7105 2.121 0.9475 ;
              RECT  1.7885 0.7105 2.121 0.753 ;
              RECT  2.0255 0.364 2.068 0.753 ;
              RECT  1.7885 0.7105 1.955 0.767 ;
              RECT  1.8735 0.3215 1.916 0.4065 ;
              RECT  1.7885 0.7105 1.831 0.9475 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.898 0.6715 0.94 0.9475 ;
              RECT  0.544 0.364 0.919 0.4065 ;
              RECT  0.8765 0.3215 0.919 0.4065 ;
              RECT  0.608 0.6715 0.94 0.714 ;
              RECT  0.622 0.364 0.6645 0.714 ;
              RECT  0.608 0.5585 0.6505 0.9475 ;
              RECT  0.544 0.3215 0.5865 0.4065 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.295 0.438 3.3515 0.7915 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.3995 0.4735 0.4985 ;
              RECT  0.265 0.544 0.4135 0.601 ;
              RECT  0.3075 0.3995 0.4135 0.601 ;
        END
    END GN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.6765 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.6765 0.042 ;
        END
    END VSS
END TLATNX4

MACRO SMDFFHQX8
    CLASS CORE ;
    SIZE 5.6565 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.4125 0.456 5.455 0.5405 ;
              RECT  4.9635 0.456 5.455 0.4985 ;
              RECT  4.974 0.4415 5.0945 0.4985 ;
              RECT  4.8505 0.491 5.006 0.5335 ;
              RECT  4.808 0.6255 4.893 0.668 ;
              RECT  4.8505 0.491 4.893 0.668 ;
        END
    END S0
    PIN D1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.077 0.569 5.342 0.6255 ;
              RECT  5.077 0.569 5.2145 0.714 ;
        END
    END D1
    PIN D0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.5395 0.6255 4.624 0.7035 ;
              RECT  4.5675 0.378 4.624 0.7035 ;
        END
    END D0
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.426 0.371 4.483 0.516 ;
              RECT  4.412 0.4595 4.4685 0.7105 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.719 0.608 3.8145 0.714 ;
              RECT  3.719 0.3995 3.7755 0.714 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.842 0.576 2.0715 0.6325 ;
              RECT  1.994 0.4525 2.0715 0.6325 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.926 0.636 0.9685 0.951 ;
              RECT  0.926 0.3745 0.9685 0.4595 ;
              RECT  0.894 0.417 0.9365 0.6785 ;
              RECT  0.636 0.523 0.9365 0.5655 ;
              RECT  0.636 0.3815 0.6785 0.951 ;
              RECT  0.042 0.424 0.6785 0.4665 ;
              RECT  0.346 0.3815 0.3885 0.951 ;
              RECT  0.0565 0.3815 0.0985 0.951 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.6565 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.6565 0.042 ;
        END
    END VSS
END SMDFFHQX8

MACRO AOI21X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.622 0.424 0.806 0.516 ;
              RECT  0.622 0.2965 0.6645 1.018 ;
              RECT  0.3955 0.2965 0.6645 0.339 ;
              RECT  0.3955 0.2545 0.438 0.339 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3955 0.24 0.7495 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.3955 0.7495 ;
              RECT  0.339 0.41 0.3955 0.7495 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.41 0.5515 0.4665 ;
              RECT  0.4665 0.41 0.523 0.735 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END AOI21X1

MACRO DFFTRX4
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.585 0.3425 4.002 0.385 ;
              RECT  3.882 0.636 3.924 0.912 ;
              RECT  3.5775 0.636 3.924 0.6785 ;
              RECT  3.5775 0.5585 3.6345 0.912 ;
              RECT  3.585 0.3425 3.6345 0.912 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.302 0.636 3.3445 0.912 ;
              RECT  2.92 0.3425 3.3375 0.385 ;
              RECT  3.012 0.636 3.3445 0.6785 ;
              RECT  3.026 0.3425 3.0685 0.6785 ;
              RECT  3.012 0.5585 3.0545 0.912 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.795 0.576 1.0145 0.6325 ;
              RECT  0.795 0.4415 1.004 0.6325 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2295 0.5585 0.3815 0.7455 ;
              RECT  0.2295 0.4875 0.286 0.7455 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.067 0.491 0.159 0.7455 ;
              RECT  0.042 0.6925 0.0985 0.7845 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END DFFTRX4

MACRO TLATNCAX3
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.298 0.714 2.3405 0.9895 ;
              RECT  2.022 0.438 2.3405 0.4805 ;
              RECT  2.298 0.3815 2.3405 0.4805 ;
              RECT  2.008 0.714 2.3405 0.7565 ;
              RECT  2.022 0.5585 2.0785 0.7565 ;
              RECT  2.022 0.3815 2.0645 0.7565 ;
              RECT  2.008 0.714 2.0505 0.9895 ;
              RECT  2.008 0.3815 2.0645 0.4665 ;
        END
    END ECK
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.548 0.576 0.6045 0.728 ;
              RECT  0.346 0.576 0.6045 0.6325 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.106 0.325 0.1625 0.5795 ;
              RECT  0.042 0.325 0.1625 0.3815 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END TLATNCAX3

MACRO FILL4
    CLASS CORE ;
    SIZE 0.5655 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.5655 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.5655 0.042 ;
        END
    END VSS
END FILL4

MACRO OAI31XL
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5935 0.6925 0.806 0.7845 ;
              RECT  0.7635 0.18 0.806 0.7845 ;
              RECT  0.5935 0.6925 0.636 0.898 ;
              RECT  0.562 0.8555 0.6045 0.94 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.424 0.0985 0.7775 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6925 0.622 ;
              RECT  0.636 0.2965 0.6925 0.622 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.431 0.523 0.7845 ;
        END
    END A2
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END OAI31XL

MACRO NOR2X1
    CLASS CORE ;
    SIZE 0.5655 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.424 0.523 0.516 ;
              RECT  0.4665 0.403 0.509 0.912 ;
              RECT  0.325 0.403 0.509 0.445 ;
              RECT  0.325 0.346 0.3675 0.445 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.403 0.24 0.7565 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.516 0.3955 0.767 ;
              RECT  0.325 0.6925 0.3815 0.8555 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.5655 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.5655 0.042 ;
        END
    END VSS
END NOR2X1

MACRO SDFFSRX4
    CLASS CORE ;
    SIZE 6.788 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.844 0.318 6.261 0.3605 ;
              RECT  6.141 0.675 6.1835 0.9225 ;
              RECT  6.109 0.608 6.1515 0.7175 ;
              RECT  5.883 0.608 6.1515 0.6505 ;
              RECT  5.883 0.5585 6.0385 0.6505 ;
              RECT  5.883 0.318 5.929 0.6505 ;
              RECT  5.851 0.647 5.9255 0.689 ;
              RECT  5.851 0.647 5.8935 0.9225 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.1795 0.318 5.5965 0.3605 ;
              RECT  5.533 0.647 5.5755 0.9225 ;
              RECT  5.243 0.647 5.5755 0.689 ;
              RECT  5.275 0.5585 5.3315 0.689 ;
              RECT  5.289 0.318 5.3315 0.689 ;
              RECT  5.243 0.647 5.2855 0.9225 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.235 0.576 3.4045 0.6325 ;
              RECT  3.235 0.392 3.2915 0.6325 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9945 0.576 3.164 0.6325 ;
              RECT  3.0475 0.392 3.104 0.6325 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0285 0.4415 1.248 0.4985 ;
              RECT  1.0285 0.4415 1.085 0.6325 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.5125 0.9475 0.714 ;
              RECT  0.8375 0.4135 0.894 0.569 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.141 0.636 0.4275 0.6925 ;
              RECT  0.141 0.569 0.258 0.6925 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7245 0.6395 0.8095 0.682 ;
              RECT  0.7245 0.1835 0.767 0.682 ;
              RECT  0.438 0.1835 0.767 0.226 ;
              RECT  0.438 0.4415 0.5405 0.4985 ;
              RECT  0.212 0.4135 0.4805 0.456 ;
              RECT  0.438 0.1835 0.4805 0.4985 ;
              RECT  0.212 0.4135 0.2545 0.4985 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.788 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.788 0.042 ;
        END
    END VSS
END SDFFSRX4

MACRO SMDFFHQX2
    CLASS CORE ;
    SIZE 4.6665 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2085 0.6185 0.251 0.926 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
              RECT  0.1975 0.3815 0.24 0.6505 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4225 0.4415 4.465 0.5265 ;
              RECT  4.267 0.4415 4.465 0.4985 ;
              RECT  4.0125 0.456 4.465 0.4985 ;
              RECT  3.8605 0.491 4.055 0.5335 ;
              RECT  3.818 0.6255 3.903 0.668 ;
              RECT  3.8605 0.491 3.903 0.668 ;
        END
    END S0
    PIN D1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.087 0.6255 4.352 0.714 ;
              RECT  4.1255 0.569 4.352 0.714 ;
        END
    END D1
    PIN D0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4965 0.601 3.6345 0.6575 ;
              RECT  3.5775 0.385 3.6345 0.6575 ;
        END
    END D0
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.369 0.4595 3.493 0.516 ;
              RECT  3.4365 0.3815 3.493 0.516 ;
              RECT  3.369 0.4595 3.4255 0.668 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.588 0.5935 2.7715 0.6505 ;
              RECT  2.715 0.4595 2.7715 0.6505 ;
              RECT  2.588 0.5585 2.6445 0.6505 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.53 0.523 0.8835 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.6665 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.6665 0.042 ;
        END
    END VSS
END SMDFFHQX2

MACRO MX4X1
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0705 0.5585 0.113 0.972 ;
              RECT  0.0565 0.2895 0.0985 0.601 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4355 0.59 2.945 0.6325 ;
              RECT  2.853 0.576 2.945 0.6325 ;
              RECT  1.7005 0.951 2.5205 0.993 ;
              RECT  2.478 0.59 2.5205 0.993 ;
              RECT  2.4355 0.59 2.5205 0.6395 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.556 0.463 2.782 0.5195 ;
              RECT  2.45 0.4415 2.662 0.4985 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.0045 0.7105 2.2165 0.767 ;
              RECT  2.04 0.569 2.0965 0.767 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7215 0.7105 1.9335 0.767 ;
              RECT  1.877 0.569 1.9335 0.767 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.3325 0.59 1.4245 0.714 ;
              RECT  1.3325 0.4415 1.389 0.714 ;
              RECT  1.2865 0.4415 1.389 0.4985 ;
        END
    END D
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.357 0.456 0.4415 0.6925 ;
              RECT  0.2825 0.4415 0.3995 0.4985 ;
        END
    END S1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END MX4X1

MACRO NOR3BX1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.318 0.424 0.3605 ;
              RECT  0.3815 0.2615 0.424 0.3605 ;
              RECT  0.173 0.8555 0.2155 0.94 ;
              RECT  0.0565 0.8555 0.2155 0.898 ;
              RECT  0.0915 0.2615 0.134 0.3605 ;
              RECT  0.0565 0.304 0.0985 0.898 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.456 0.6645 0.8095 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.24 0.7845 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END NOR3BX1

MACRO SDFFX1
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.516 ;
              RECT  0.608 0.3815 0.6505 0.9295 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.141 0.3815 0.1975 0.912 ;
              RECT  0.042 0.424 0.1975 0.516 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.486 0.4415 3.652 0.4985 ;
              RECT  3.486 0.4135 3.528 0.4985 ;
              RECT  3.097 0.4525 3.652 0.4945 ;
              RECT  3.0545 0.6395 3.1395 0.682 ;
              RECT  3.097 0.4525 3.1395 0.682 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.3655 0.6045 3.684 0.661 ;
              RECT  3.4185 0.569 3.684 0.661 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.814 0.4595 2.8705 0.682 ;
              RECT  2.729 0.4595 2.8705 0.516 ;
              RECT  2.729 0.4135 2.786 0.516 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8485 0.53 0.905 0.6785 ;
              RECT  0.7315 0.7105 0.898 0.767 ;
              RECT  0.841 0.622 0.898 0.767 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END SDFFX1

MACRO AND2X6
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.354 0.636 1.3965 0.9685 ;
              RECT  0.7635 0.371 1.3855 0.4135 ;
              RECT  1.3435 0.194 1.3855 0.4135 ;
              RECT  0.774 0.636 1.3965 0.6785 ;
              RECT  1.1735 0.5585 1.23 0.6785 ;
              RECT  1.1735 0.371 1.216 0.6785 ;
              RECT  1.064 0.636 1.1065 0.9685 ;
              RECT  1.0535 0.194 1.096 0.4135 ;
              RECT  0.774 0.636 0.8165 0.9685 ;
              RECT  0.7635 0.194 0.806 0.4135 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2015 0.555 0.4665 0.6115 ;
              RECT  0.2015 0.555 0.3995 0.7 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.537 0.4415 0.5795 0.5335 ;
              RECT  0.0245 0.4415 0.5795 0.484 ;
              RECT  0.088 0.4415 0.1305 0.5515 ;
              RECT  0.0245 0.4415 0.1305 0.5055 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END AND2X6

MACRO SEDFFHQX8
    CLASS CORE ;
    SIZE 6.2225 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  6.0455 0.456 6.088 0.5405 ;
              RECT  5.6815 0.456 6.088 0.4985 ;
              RECT  5.487 0.449 5.7735 0.491 ;
              RECT  5.6815 0.4415 5.7735 0.4985 ;
              RECT  5.487 0.449 5.5295 0.714 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.918 0.569 5.975 0.76 ;
              RECT  5.7555 0.569 5.975 0.6325 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.1335 0.438 5.19 0.7915 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.3025 0.4525 4.458 0.509 ;
              RECT  4.267 0.576 4.359 0.6715 ;
              RECT  4.3025 0.4525 4.359 0.6715 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8805 0.4945 1.937 0.795 ;
              RECT  1.8275 0.4945 1.937 0.6505 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.926 0.636 0.9685 0.951 ;
              RECT  0.926 0.371 0.9685 0.456 ;
              RECT  0.894 0.4135 0.9365 0.6785 ;
              RECT  0.346 0.523 0.9365 0.5655 ;
              RECT  0.636 0.3815 0.6785 0.951 ;
              RECT  0.346 0.3815 0.3885 0.951 ;
              RECT  0.042 0.456 0.3885 0.4985 ;
              RECT  0.0565 0.3815 0.0985 0.951 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.2225 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.2225 0.042 ;
        END
    END VSS
END SEDFFHQX8

MACRO DFFTRX2
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.892 0.403 3.005 0.4595 ;
              RECT  2.906 0.622 2.9625 0.912 ;
              RECT  2.892 0.403 2.9485 0.6645 ;
              RECT  2.8705 0.424 2.9485 0.516 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.63 0.403 2.6725 0.912 ;
              RECT  2.588 0.403 2.6725 0.516 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.2485 0.544 2.404 0.6325 ;
              RECT  2.305 0.378 2.3615 0.6325 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0845 0.4065 0.141 0.7175 ;
              RECT  0.042 0.4065 0.141 0.516 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END DFFTRX2

MACRO TLATNTSCAX4
    CLASS CORE ;
    SIZE 2.9695 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4065 0.7105 0.576 0.8305 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.576 0.654 0.6395 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.067 0.484 0.1235 0.7495 ;
              RECT  0.042 0.6925 0.0985 0.813 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7255 0.3285 2.768 0.979 ;
              RECT  2.4465 0.4735 2.768 0.516 ;
              RECT  2.4675 0.4735 2.51 0.728 ;
              RECT  2.4465 0.424 2.503 0.516 ;
              RECT  2.4465 0.3285 2.489 0.516 ;
              RECT  2.4355 0.6855 2.478 0.979 ;
              RECT  2.4355 0.3285 2.489 0.4135 ;
        END
    END ECK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.9695 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.9695 0.042 ;
        END
    END VSS
END TLATNTSCAX4

MACRO DFFQX4
    CLASS CORE ;
    SIZE 2.9695 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.464 0.576 2.662 0.6325 ;
              RECT  2.464 0.477 2.5205 0.689 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.325 0.24 0.6785 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7385 0.3425 0.8375 0.385 ;
              RECT  0.7565 0.682 0.799 0.958 ;
              RECT  0.7385 0.3425 0.781 0.721 ;
              RECT  0.4665 0.4735 0.781 0.516 ;
              RECT  0.4665 0.424 0.523 0.516 ;
              RECT  0.4665 0.3425 0.509 0.958 ;
              RECT  0.4205 0.3425 0.509 0.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.9695 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.9695 0.042 ;
        END
    END VSS
END DFFQX4

MACRO AND3X8
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.983 0.403 2.0785 0.445 ;
              RECT  2.015 0.6575 2.0575 0.972 ;
              RECT  1.177 0.4135 2.015 0.456 ;
              RECT  1.1455 0.6575 2.0575 0.7 ;
              RECT  1.8805 0.4135 1.937 0.516 ;
              RECT  1.8805 0.4135 1.923 0.7 ;
              RECT  1.704 0.403 1.7885 0.456 ;
              RECT  1.725 0.6575 1.7675 0.972 ;
              RECT  1.414 0.403 1.499 0.456 ;
              RECT  1.435 0.6575 1.4775 0.972 ;
              RECT  1.124 0.403 1.209 0.445 ;
              RECT  1.1455 0.6575 1.1875 0.972 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.445 0.576 0.608 0.7035 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.463 0.806 0.6505 ;
              RECT  0.41 0.463 0.806 0.5055 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.898 0.35 0.94 0.5195 ;
              RECT  0.1975 0.35 0.94 0.392 ;
              RECT  0.1835 0.424 0.24 0.537 ;
              RECT  0.1975 0.35 0.24 0.537 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END AND3X8

MACRO AOI221X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0465 0.1555 1.0885 1.032 ;
              RECT  0.615 0.2965 1.0885 0.339 ;
              RECT  1.032 0.1555 1.0885 0.339 ;
              RECT  0.5655 0.2825 0.6505 0.325 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.41 0.6645 0.7635 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.41 0.806 0.7635 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.318 0.24 0.6715 ;
        END
    END A0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.4595 0.9755 0.516 ;
              RECT  0.8905 0.41 0.9475 0.735 ;
        END
    END C0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.1555 0.3815 0.509 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END AOI221X1

MACRO TLATNX2
    CLASS CORE ;
    SIZE 2.5455 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.5455 0.042 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.5455 1.209 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.484 0.3995 0.5405 ;
              RECT  0.1375 0.576 0.364 0.6325 ;
              RECT  0.3075 0.484 0.364 0.6325 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.29 0.4415 1.3965 0.6325 ;
        END
    END GN
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.325 1.6545 0.912 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1955 0.4415 2.379 0.4985 ;
              RECT  2.1955 0.325 2.252 0.912 ;
        END
    END Q
END TLATNX2

MACRO INVXL
    CLASS CORE ;
    SIZE 0.2825 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2085 0.636 0.265 0.6925 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.509 0.1375 0.5655 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.2825 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.2825 0.042 ;
        END
    END VSS
END INVXL

MACRO ADDFXL
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.729 0.424 2.786 0.516 ;
              RECT  2.729 0.2085 2.7715 0.8485 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2225 0.608 0.265 0.7385 ;
              RECT  0.0565 0.339 0.265 0.3815 ;
              RECT  0.2225 0.2015 0.265 0.3815 ;
              RECT  0.042 0.608 0.265 0.6505 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
              RECT  0.0565 0.339 0.0985 0.6505 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.393 0.5795 2.3755 0.622 ;
              RECT  0.7455 0.5975 1.435 0.6395 ;
              RECT  1.117 0.5975 1.248 0.767 ;
              RECT  0.7455 0.555 0.788 0.6395 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4465 0.4665 2.503 0.7105 ;
              RECT  0.9435 0.4665 2.503 0.509 ;
              RECT  0.6325 0.456 0.986 0.484 ;
              RECT  0.8375 0.4665 2.503 0.4985 ;
              RECT  0.6325 0.4415 0.873 0.484 ;
              RECT  0.5865 0.4735 0.675 0.516 ;
        END
    END A
    PIN CI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.057 0.3535 2.227 0.3955 ;
              RECT  1.057 0.3075 1.248 0.3955 ;
        END
    END CI
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END ADDFXL

MACRO INVX6
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.76 0.4945 0.8165 0.5655 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.509 0.106 0.615 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END INVX6

MACRO XNOR3XL
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.998 0.735 3.0865 0.7775 ;
              RECT  3.044 0.403 3.0865 0.7775 ;
              RECT  2.9945 0.4415 3.0865 0.4985 ;
              RECT  2.998 0.403 3.0865 0.4985 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.067 0.449 0.1235 0.7775 ;
              RECT  0.042 0.5585 0.1235 0.6505 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.4945 0.3815 0.7775 ;
              RECT  0.3075 0.4415 0.364 0.5515 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.146 0.6185 2.379 0.661 ;
              RECT  2.146 0.576 2.2375 0.661 ;
              RECT  2.146 0.47 2.188 0.661 ;
              RECT  2.068 0.47 2.188 0.5125 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END XNOR3XL

MACRO OR4X2
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.2825 1.23 0.958 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5935 0.339 0.6505 0.53 ;
              RECT  0.4665 0.424 0.6505 0.4805 ;
              RECT  0.4665 0.424 0.523 0.516 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5585 0.3955 0.6785 ;
              RECT  0.339 0.339 0.3955 0.6785 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5585 0.2545 0.6785 ;
              RECT  0.1975 0.339 0.2545 0.6785 ;
        END
    END D
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8445 0.4415 0.965 0.4985 ;
              RECT  0.8445 0.247 0.9015 0.537 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END OR4X2

MACRO AO21X1
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8625 0.339 0.905 1.0465 ;
              RECT  0.7495 0.339 0.905 0.3815 ;
              RECT  0.7495 0.2895 0.806 0.3815 ;
              RECT  0.7635 0.2615 0.806 0.3815 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.318 0.24 0.6715 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.1555 0.3815 0.509 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5585 0.523 0.7775 ;
              RECT  0.4595 0.431 0.516 0.643 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END AO21X1

MACRO OAI221XL
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.103 0.827 1.23 0.919 ;
              RECT  0.654 0.788 1.2055 0.8305 ;
              RECT  1.163 0.2295 1.2055 0.919 ;
              RECT  0.654 0.788 0.6965 0.919 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.477 0.24 0.8305 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.456 0.576 0.8095 0.6325 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3285 0.569 0.385 0.8835 ;
              RECT  0.325 0.827 0.3815 0.919 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.364 0.9475 0.7175 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.3675 1.092 0.7175 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OAI221XL

MACRO NOR3X1
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.5585 0.6645 0.6505 ;
              RECT  0.608 0.346 0.6505 0.912 ;
              RECT  0.318 0.403 0.6505 0.445 ;
              RECT  0.318 0.247 0.3605 0.445 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4805 0.516 0.537 0.7845 ;
              RECT  0.4665 0.6925 0.523 0.8555 ;
        END
    END C
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.403 0.24 0.7565 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.516 0.3815 0.8695 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END NOR3X1

MACRO AND2X4
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.424 1.0885 0.516 ;
              RECT  0.689 0.7705 1.0745 0.813 ;
              RECT  1.032 0.311 1.0745 0.813 ;
              RECT  0.9895 0.7705 1.032 1.0465 ;
              RECT  0.9895 0.2685 1.032 0.3535 ;
              RECT  0.7175 0.311 1.0745 0.3535 ;
              RECT  0.668 0.2965 0.753 0.339 ;
              RECT  0.689 0.7705 0.7315 1.0465 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.537 0.523 0.8905 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.226 0.4415 0.2825 0.576 ;
              RECT  0.042 0.4415 0.2825 0.4985 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END AND2X4

MACRO TLATNCAX12
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.431 0.6575 1.6545 0.7 ;
              RECT  0.431 0.3605 1.633 0.403 ;
              RECT  1.5905 0.1835 1.633 0.403 ;
              RECT  1.301 0.1835 1.3435 0.403 ;
              RECT  1.011 0.1835 1.0535 0.403 ;
              RECT  0.431 0.636 0.806 0.7 ;
              RECT  0.7 0.5585 0.806 0.7 ;
              RECT  0.721 0.1835 0.7635 0.403 ;
              RECT  0.7 0.3605 0.742 0.7 ;
              RECT  0.431 0.636 0.4735 0.721 ;
              RECT  0.431 0.1835 0.4735 0.403 ;
        END
    END ECK
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.719 0.6925 3.7755 0.8625 ;
              RECT  3.627 0.6925 3.7755 0.7495 ;
              RECT  3.627 0.601 3.684 0.7495 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.576 0.3605 0.6325 ;
              RECT  0.166 0.438 0.2295 0.6325 ;
              RECT  0.1445 0.438 0.2295 0.4945 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END TLATNCAX12

MACRO XOR2X4
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.951 0.5265 1.0355 ;
              RECT  0.484 0.233 0.5265 0.318 ;
              RECT  0.4525 0.76 0.4945 0.993 ;
              RECT  0.1835 0.3885 0.4945 0.431 ;
              RECT  0.4525 0.2755 0.4945 0.431 ;
              RECT  0.1835 0.76 0.4945 0.8025 ;
              RECT  0.173 0.3535 0.258 0.3955 ;
              RECT  0.1835 0.6925 0.24 0.8025 ;
              RECT  0.1835 0.6925 0.2365 1.0355 ;
              RECT  0.1835 0.3535 0.226 1.0355 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5025 0.4415 1.559 0.5265 ;
              RECT  1.2335 0.4415 1.559 0.4985 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6785 0.502 0.8235 0.767 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END XOR2X4

MACRO SDFFSX1
    CLASS CORE ;
    SIZE 4.9495 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8445 0.3815 0.887 0.735 ;
              RECT  0.7635 0.636 0.887 0.735 ;
              RECT  0.7635 0.636 0.806 0.912 ;
              RECT  0.7495 0.6925 0.806 0.7845 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.403 0.3815 0.6925 ;
              RECT  0.2965 0.636 0.3535 0.912 ;
              RECT  0.2755 0.403 0.3815 0.4595 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.7125 0.4135 4.755 0.4985 ;
              RECT  4.4935 0.456 4.755 0.4985 ;
              RECT  4.4935 0.4415 4.642 0.4985 ;
              RECT  4.2955 0.463 4.5925 0.5055 ;
              RECT  4.4935 0.4135 4.536 0.5055 ;
              RECT  4.253 0.615 4.338 0.6575 ;
              RECT  4.2955 0.463 4.338 0.6575 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.5675 0.576 4.734 0.661 ;
              RECT  4.4085 0.576 4.734 0.6325 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.8605 0.509 4.069 0.5655 ;
              RECT  3.8605 0.364 3.917 0.5655 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.7335 0.364 3.79 0.7035 ;
              RECT  3.719 0.3885 3.79 0.516 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4005 0.233 2.485 0.2755 ;
              RECT  2.1315 0.247 2.443 0.2895 ;
              RECT  1.58 0.2295 2.174 0.272 ;
              RECT  1.3115 0.59 1.672 0.6325 ;
              RECT  1.58 0.576 1.672 0.6325 ;
              RECT  1.58 0.2295 1.6225 0.6325 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.9495 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.9495 0.042 ;
        END
    END VSS
END SDFFSX1

MACRO AOI2BB2X4
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.754 0.7035 2.7965 0.788 ;
              RECT  1.863 0.7035 2.7965 0.7455 ;
              RECT  2.6335 0.3145 2.676 0.7455 ;
              RECT  2.588 0.3145 2.676 0.357 ;
              RECT  2.464 0.7035 2.5065 0.788 ;
              RECT  2.174 0.7035 2.2165 0.788 ;
              RECT  1.8735 0.3145 2.114 0.357 ;
              RECT  1.884 0.7035 1.955 0.788 ;
              RECT  1.039 0.3285 1.909 0.371 ;
              RECT  1.863 0.569 1.9055 0.767 ;
              RECT  1.75 0.569 1.9055 0.6115 ;
              RECT  1.75 0.3285 1.7925 0.6115 ;
              RECT  1.428 0.3145 1.513 0.371 ;
              RECT  0.9895 0.3145 1.0745 0.357 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1 0.576 2.563 0.6325 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.747 0.4525 2.8705 0.4945 ;
              RECT  2.747 0.2015 2.7895 0.4945 ;
              RECT  2.4745 0.2015 2.7895 0.2435 ;
              RECT  1.863 0.456 2.517 0.4985 ;
              RECT  2.4745 0.2015 2.517 0.4985 ;
              RECT  1.863 0.4415 1.955 0.4985 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.491 0.3815 0.8445 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.491 0.24 0.8445 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END AOI2BB2X4

MACRO NOR4BX1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6855 0.24 0.728 0.325 ;
              RECT  0.0565 0.318 0.6925 0.3605 ;
              RECT  0.6505 0.2825 0.728 0.325 ;
              RECT  0.385 0.2615 0.4275 0.3605 ;
              RECT  0.311 0.8555 0.3535 1.0075 ;
              RECT  0.0565 0.8555 0.3535 0.898 ;
              RECT  0.0565 0.318 0.0985 0.898 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.431 1.0885 0.7845 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7315 0.5725 0.9615 0.6325 ;
              RECT  0.6115 0.5725 0.9615 0.629 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.449 0.449 0.5405 0.767 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.24 0.7845 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END NOR4BX1

MACRO SEDFFTRX1
    CLASS CORE ;
    SIZE 5.798 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.8325 0.424 3.917 0.516 ;
              RECT  3.758 0.707 3.889 0.7635 ;
              RECT  3.8325 0.3815 3.889 0.7635 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.3815 0.0985 0.912 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.579 0.4945 5.6355 0.7495 ;
              RECT  5.5575 0.6925 5.614 0.827 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.275 0.544 5.3315 0.6505 ;
              RECT  4.939 0.544 5.3315 0.601 ;
        END
    END E
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1435 0.6185 4.32 0.675 ;
              RECT  4.1435 0.6185 4.2 0.852 ;
        END
    END RN
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8845 0.4525 3.0685 0.6505 ;
              RECT  2.8845 0.4525 2.9415 0.6785 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.2525 0.339 3.295 0.5795 ;
              RECT  2.7715 0.339 3.295 0.3815 ;
              RECT  2.7715 0.339 2.814 0.5795 ;
              RECT  2.7115 0.4415 2.814 0.4985 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.4735 2.3685 0.7915 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.798 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.798 0.042 ;
        END
    END VSS
END SEDFFTRX1

MACRO SEDFFTRX4
    CLASS CORE ;
    SIZE 6.788 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1255 0.346 4.543 0.3885 ;
              RECT  4.32 0.7245 4.451 0.767 ;
              RECT  4.1255 0.7105 4.3625 0.753 ;
              RECT  4.034 0.7245 4.2175 0.767 ;
              RECT  4.175 0.346 4.2175 0.767 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.461 0.325 3.878 0.3675 ;
              RECT  3.7225 0.7105 3.765 0.795 ;
              RECT  3.56 0.7105 3.765 0.753 ;
              RECT  3.348 0.7245 3.652 0.767 ;
              RECT  3.5775 0.325 3.62 0.767 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  6.5475 0.2895 6.604 0.643 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.9605 0.5935 6.3285 0.6505 ;
              RECT  6.272 0.523 6.3285 0.6505 ;
              RECT  6.2645 0.5585 6.3285 0.6505 ;
        END
    END E
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.1335 0.5515 5.2255 0.8695 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.424 3.21 0.735 ;
              RECT  3.111 0.4595 3.21 0.516 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.134 0.6395 0.417 0.6965 ;
              RECT  0.134 0.569 0.41 0.6965 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.714 0.212 0.7565 0.601 ;
              RECT  0.385 0.212 0.7565 0.2545 ;
              RECT  0.159 0.456 0.53 0.4985 ;
              RECT  0.385 0.212 0.4275 0.4985 ;
              RECT  0.159 0.4415 0.258 0.4985 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.788 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.788 0.042 ;
        END
    END VSS
END SEDFFTRX4

MACRO NAND3BX1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.392 0.8485 0.4345 1.0465 ;
              RECT  0.042 0.8485 0.4345 0.8905 ;
              RECT  0.0565 0.311 0.1835 0.3535 ;
              RECT  0.141 0.2685 0.1835 0.3535 ;
              RECT  0.1025 0.8485 0.1445 1.0465 ;
              RECT  0.042 0.6925 0.0985 0.8905 ;
              RECT  0.0565 0.311 0.0985 0.8905 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.537 0.6645 0.8905 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.424 0.3815 0.7775 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END NAND3BX1

MACRO DFFQX2
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1775 0.3815 2.22 0.6505 ;
              RECT  2.1635 0.5585 2.206 0.958 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.689 0.4595 0.7455 0.689 ;
              RECT  0.608 0.4595 0.7455 0.516 ;
              RECT  0.608 0.417 0.6645 0.516 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.205 0.4415 0.2615 0.615 ;
              RECT  0.042 0.4415 0.2615 0.516 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END DFFQX2

MACRO AND3X6
    CLASS CORE ;
    SIZE 1.838 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.711 0.6505 1.7535 0.9685 ;
              RECT  1.131 0.4205 1.7535 0.463 ;
              RECT  1.711 0.2435 1.7535 0.463 ;
              RECT  1.131 0.6505 1.7535 0.6925 ;
              RECT  1.598 0.5585 1.6545 0.6925 ;
              RECT  1.598 0.4205 1.64 0.6925 ;
              RECT  1.421 0.6505 1.4635 0.9685 ;
              RECT  1.421 0.2435 1.4635 0.463 ;
              RECT  1.131 0.6505 1.1735 0.9685 ;
              RECT  1.131 0.2435 1.1735 0.463 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3745 0.576 0.6785 0.682 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.463 0.806 0.6505 ;
              RECT  0.332 0.463 0.806 0.5055 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.35 0.933 0.53 ;
              RECT  0.219 0.35 0.933 0.392 ;
              RECT  0.219 0.35 0.2615 0.5195 ;
              RECT  0.1835 0.424 0.2615 0.516 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.838 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.838 0.042 ;
        END
    END VSS
END AND3X6

MACRO AOI221X4
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.0015 0.7035 3.044 0.8025 ;
              RECT  1.347 0.7035 3.044 0.7455 ;
              RECT  2.9095 0.3145 2.9945 0.357 ;
              RECT  0.5865 0.3285 2.945 0.371 ;
              RECT  2.7115 0.7035 2.754 0.8025 ;
              RECT  2.5985 0.3145 2.683 0.371 ;
              RECT  2.2165 0.3145 2.3015 0.371 ;
              RECT  1.6755 0.3145 1.7605 0.371 ;
              RECT  1.347 0.3285 1.389 0.7455 ;
              RECT  1.2975 0.4415 1.389 0.4985 ;
              RECT  0.9755 0.3145 1.0605 0.371 ;
              RECT  0.537 0.3145 0.622 0.357 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.576 1.0075 0.6325 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7675 0.576 2.2485 0.6325 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1625 0.456 1.2265 0.4985 ;
              RECT  0.166 0.4415 0.258 0.4985 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4215 0.576 2.5205 0.6325 ;
              RECT  1.4775 0.463 2.5065 0.5055 ;
              RECT  2.4215 0.463 2.464 0.6325 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7115 0.445 2.966 0.502 ;
              RECT  2.7115 0.4415 2.8035 0.6325 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END AOI221X4

MACRO XOR2X2
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.265 0.8165 0.3075 0.9015 ;
              RECT  0.1975 0.35 0.3075 0.392 ;
              RECT  0.265 0.3075 0.3075 0.392 ;
              RECT  0.1975 0.8165 0.3075 0.859 ;
              RECT  0.1975 0.35 0.24 0.859 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9435 0.576 1.262 0.6185 ;
              RECT  1.0145 0.576 1.1065 0.6325 ;
              RECT  0.7495 0.583 1.1065 0.6255 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.509 0.576 0.5655 0.8445 ;
              RECT  0.424 0.576 0.5655 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END XOR2X2

MACRO DFFRX4
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.581 0.403 3.9985 0.445 ;
              RECT  3.864 0.753 3.9065 0.94 ;
              RECT  3.574 0.742 3.882 0.7845 ;
              RECT  3.8395 0.753 3.9065 0.799 ;
              RECT  3.5775 0.6925 3.6345 0.7845 ;
              RECT  3.581 0.403 3.6345 0.7845 ;
              RECT  3.574 0.742 3.6165 0.94 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9165 0.3885 3.334 0.431 ;
              RECT  3.27 0.6645 3.3125 0.94 ;
              RECT  2.98 0.6645 3.3125 0.707 ;
              RECT  3.012 0.5585 3.0685 0.707 ;
              RECT  3.012 0.3885 3.0545 0.707 ;
              RECT  2.98 0.6645 3.0225 0.94 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3405 0.403 2.761 0.445 ;
              RECT  2.3405 0.2895 2.3825 0.445 ;
              RECT  2.135 0.2895 2.3825 0.332 ;
              RECT  2.135 0.212 2.1775 0.332 ;
              RECT  1.6545 0.212 2.1775 0.2545 ;
              RECT  1.3045 0.5725 1.697 0.615 ;
              RECT  1.6545 0.212 1.697 0.615 ;
              RECT  1.58 0.4415 1.697 0.4985 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.555 0.7245 0.6115 ;
              RECT  0.608 0.555 0.6645 0.8485 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.1765 0.615 ;
              RECT  0.12 0.3745 0.1765 0.615 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END DFFRX4

MACRO AND4X8
    CLASS CORE ;
    SIZE 2.5455 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4355 0.636 2.478 0.951 ;
              RECT  1.566 0.636 2.478 0.6785 ;
              RECT  2.319 0.339 2.4145 0.3815 ;
              RECT  1.513 0.35 2.3615 0.392 ;
              RECT  2.1635 0.5585 2.22 0.6785 ;
              RECT  2.1635 0.35 2.206 0.6785 ;
              RECT  2.146 0.636 2.188 0.951 ;
              RECT  2.04 0.339 2.1245 0.392 ;
              RECT  1.856 0.636 1.8985 0.951 ;
              RECT  1.75 0.339 1.8345 0.392 ;
              RECT  1.566 0.636 1.6085 0.951 ;
              RECT  1.46 0.339 1.5555 0.3815 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.795 1.276 0.8375 ;
              RECT  1.2335 0.5795 1.276 0.8375 ;
              RECT  1.1735 0.6925 1.276 0.8375 ;
              RECT  0.1835 0.5795 0.226 0.8375 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0605 0.537 1.163 0.622 ;
              RECT  0.325 0.682 1.103 0.7245 ;
              RECT  1.0605 0.537 1.103 0.7245 ;
              RECT  0.325 0.5585 0.3815 0.7245 ;
              RECT  0.2965 0.59 0.3815 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4735 0.569 0.9755 0.6115 ;
              RECT  0.933 0.4415 0.9755 0.6115 ;
              RECT  0.873 0.4415 0.9755 0.4985 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.4415 0.8025 0.4985 ;
              RECT  0.608 0.2825 0.6645 0.4985 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.5455 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.5455 0.042 ;
        END
    END VSS
END AND4X8

MACRO SDFFRXL
    CLASS CORE ;
    SIZE 4.2425 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.6925 0.6645 0.979 ;
              RECT  0.608 0.332 0.6505 0.979 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1445 0.3815 0.2015 0.721 ;
              RECT  0.042 0.424 0.2015 0.516 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.9845 0.4415 4.076 0.4985 ;
              RECT  3.9845 0.3285 4.0265 0.4985 ;
              RECT  3.3975 0.3285 4.0265 0.371 ;
              RECT  3.585 0.3285 3.627 0.5125 ;
              RECT  3.3975 0.3285 3.44 0.643 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.698 0.5795 3.9135 0.636 ;
              RECT  3.698 0.4415 3.7935 0.636 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.157 0.35 3.2135 0.615 ;
              RECT  3.1535 0.5585 3.21 0.7 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.5795 1.4915 0.636 ;
              RECT  1.156 0.576 1.248 0.6505 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.799 0.5865 0.8555 0.767 ;
              RECT  0.7495 0.6925 0.806 0.8905 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.2425 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.2425 0.042 ;
        END
    END VSS
END SDFFRXL

MACRO SDFFNSRX1
    CLASS CORE ;
    SIZE 5.515 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6645 0.364 0.707 0.449 ;
              RECT  0.661 0.7315 0.7035 1.0075 ;
              RECT  0.608 0.6925 0.6715 0.7845 ;
              RECT  0.629 0.392 0.6715 0.7845 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.912 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.978 0.456 5.317 0.5125 ;
              RECT  5.1155 0.4415 5.2075 0.5125 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.091 0.583 5.317 0.767 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.5675 0.6925 4.6385 0.813 ;
              RECT  4.582 0.4735 4.6385 0.813 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4405 0.4735 4.497 0.813 ;
              RECT  4.426 0.4735 4.497 0.6505 ;
        END
    END CKN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8705 0.951 3.1925 0.993 ;
              RECT  2.8705 0.8305 2.913 0.993 ;
              RECT  2.234 0.8305 2.913 0.873 ;
              RECT  2.234 0.654 2.2765 0.873 ;
              RECT  1.6295 0.654 2.2765 0.6965 ;
              RECT  1.6295 0.576 1.672 0.6965 ;
              RECT  1.506 0.59 1.672 0.6325 ;
              RECT  1.58 0.576 1.672 0.6325 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.774 0.7105 0.965 0.852 ;
              RECT  0.88 0.6325 0.965 0.852 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.515 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.515 0.042 ;
        END
    END VSS
END SDFFNSRX1

MACRO AOI31X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.424 0.806 0.516 ;
              RECT  0.7495 0.318 0.7915 1.0465 ;
              RECT  0.516 0.318 0.7915 0.3605 ;
              RECT  0.516 0.2615 0.5585 0.3605 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.318 0.24 0.6715 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.431 0.6645 0.7845 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4595 0.431 0.523 0.6505 ;
              RECT  0.4595 0.431 0.516 0.7775 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.332 0.1905 0.3885 0.502 ;
              RECT  0.325 0.1555 0.3815 0.247 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END AOI31X1

MACRO SDFFNSRX4
    CLASS CORE ;
    SIZE 6.6465 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.713 0.339 6.1305 0.3815 ;
              RECT  5.9785 0.647 6.021 0.9225 ;
              RECT  5.6885 0.647 6.021 0.689 ;
              RECT  5.699 0.5585 5.7555 0.689 ;
              RECT  5.713 0.339 5.7555 0.689 ;
              RECT  5.6885 0.647 5.731 0.9225 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.0485 0.339 5.4655 0.3815 ;
              RECT  5.3985 0.608 5.441 0.9225 ;
              RECT  5.1335 0.608 5.441 0.6505 ;
              RECT  5.1335 0.5585 5.19 0.6505 ;
              RECT  5.1085 0.647 5.176 0.9225 ;
              RECT  5.1335 0.339 5.176 0.9225 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8885 0.463 3.2455 0.5195 ;
              RECT  2.853 0.4415 2.945 0.4985 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7255 0.4415 2.782 0.6395 ;
              RECT  2.57 0.4415 2.782 0.4985 ;
        END
    END SN
    PIN CKN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.4945 1.0885 0.8485 ;
        END
    END CKN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.4595 0.9475 0.813 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.5055 0.4805 0.6505 ;
              RECT  0.325 0.5055 0.3815 0.76 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7775 0.2085 0.82 0.7495 ;
              RECT  0.5515 0.2085 0.82 0.251 ;
              RECT  0.5515 0.2085 0.5935 0.562 ;
              RECT  0.212 0.392 0.5935 0.4345 ;
              RECT  0.4665 0.2895 0.5935 0.4345 ;
              RECT  0.212 0.392 0.2545 0.477 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.6465 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.6465 0.042 ;
        END
    END VSS
END SDFFNSRX4

MACRO AND2X2
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.516 ;
              RECT  0.608 0.3145 0.6505 0.9475 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3605 0.484 0.417 0.8025 ;
              RECT  0.325 0.484 0.417 0.6505 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0845 0.484 0.141 0.7845 ;
              RECT  0.042 0.675 0.0985 0.795 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END AND2X2

MACRO OR3XL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.622 0.728 0.806 0.7845 ;
              RECT  0.7495 0.1835 0.806 0.7845 ;
              RECT  0.622 0.728 0.6785 0.8555 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4415 0.7105 0.5405 0.767 ;
              RECT  0.4415 0.456 0.4985 0.767 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2015 0.4525 0.258 0.788 ;
              RECT  0.1835 0.4525 0.258 0.6505 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.4345 0.0985 0.788 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OR3XL

MACRO CLKBUFX4
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4735 0.2825 0.5585 0.325 ;
              RECT  0.4945 0.6925 0.537 0.9685 ;
              RECT  0.1625 0.2965 0.509 0.339 ;
              RECT  0.1625 0.6925 0.537 0.735 ;
              RECT  0.1835 0.6925 0.24 0.7845 ;
              RECT  0.1835 0.6925 0.2365 0.9685 ;
              RECT  0.194 0.2545 0.2365 0.339 ;
              RECT  0.1625 0.2965 0.205 0.735 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.5515 0.728 0.608 ;
              RECT  0.6715 0.523 0.728 0.608 ;
              RECT  0.608 0.5515 0.6645 0.813 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END CLKBUFX4

MACRO AO22X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0885 0.742 1.131 1.018 ;
              RECT  1.032 0.6925 1.0885 0.7845 ;
              RECT  1.032 0.293 1.0745 0.7845 ;
              RECT  1.0285 0.293 1.0745 0.378 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7245 0.5585 0.806 0.707 ;
              RECT  0.7245 0.463 0.781 0.7915 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.445 0.113 0.7495 ;
              RECT  0.042 0.6925 0.0985 0.7845 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.449 0.4415 0.5405 0.5265 ;
              RECT  0.449 0.4415 0.5055 0.76 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3215 0.5585 0.378 0.7385 ;
              RECT  0.1835 0.5585 0.378 0.615 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END AO22X1

MACRO NOR4X1
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.403 0.9475 0.516 ;
              RECT  0.8765 0.403 0.919 0.912 ;
              RECT  0.403 0.403 0.9475 0.445 ;
              RECT  0.7 0.346 0.742 0.445 ;
              RECT  0.403 0.346 0.445 0.445 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2755 0.424 0.332 0.5515 ;
              RECT  0.042 0.424 0.332 0.4805 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4805 0.516 0.537 0.7495 ;
              RECT  0.4665 0.6925 0.523 0.8555 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.516 0.6645 0.8695 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.516 0.806 0.8695 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END NOR4X1

MACRO NAND3BX4
    CLASS CORE ;
    SIZE 2.121 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.6615 0.795 1.704 1.0075 ;
              RECT  0.212 0.795 1.704 0.8375 ;
              RECT  1.3715 0.795 1.414 1.0075 ;
              RECT  0.042 0.2895 1.3785 0.332 ;
              RECT  1.0815 0.795 1.124 1.0075 ;
              RECT  0.7915 0.795 0.834 1.0075 ;
              RECT  0.502 0.795 0.544 1.0075 ;
              RECT  0.212 0.7315 0.2545 1.0075 ;
              RECT  0.0565 0.7315 0.2545 0.774 ;
              RECT  0.0565 0.2895 0.0985 0.774 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1345 0.569 1.6015 0.6115 ;
              RECT  0.866 0.5265 1.177 0.569 ;
              RECT  0.4665 0.569 0.9085 0.6115 ;
              RECT  0.4665 0.463 0.509 0.6115 ;
              RECT  0.2825 0.463 0.509 0.5055 ;
              RECT  0.3075 0.4415 0.3995 0.5055 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.757 0.5055 1.962 0.562 ;
              RECT  1.757 0.4415 1.8135 0.562 ;
              RECT  1.672 0.4415 1.8135 0.4985 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.248 0.456 1.3325 0.4985 ;
              RECT  0.753 0.4135 1.29 0.456 ;
              RECT  0.5795 0.456 0.795 0.4985 ;
              RECT  0.59 0.4415 0.682 0.4985 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.121 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.121 0.042 ;
        END
    END VSS
END NAND3BX4

MACRO AND3X4
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0355 0.5585 1.23 0.6505 ;
              RECT  0.735 0.7635 1.078 0.806 ;
              RECT  1.0355 0.403 1.078 0.806 ;
              RECT  1.025 0.7635 1.0675 1.039 ;
              RECT  0.682 0.417 1.078 0.4595 ;
              RECT  0.9435 0.403 1.078 0.4595 ;
              RECT  0.735 0.7635 0.7775 1.039 ;
              RECT  0.6325 0.403 0.7175 0.445 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.6925 0.6645 0.8835 ;
              RECT  0.4945 0.6925 0.6645 0.7495 ;
              RECT  0.4945 0.643 0.5515 0.7495 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2545 0.4595 0.311 0.707 ;
              RECT  0.1835 0.4595 0.311 0.516 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.417 0.0985 0.7705 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END AND3X4

MACRO DFFRHQX1
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1025 0.647 0.159 0.9225 ;
              RECT  0.0635 0.272 0.12 0.357 ;
              RECT  0.042 0.647 0.159 0.7035 ;
              RECT  0.042 0.3075 0.0985 0.7035 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9755 0.6505 1.248 0.714 ;
              RECT  1.156 0.576 1.248 0.714 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3425 0.5265 0.4525 0.583 ;
              RECT  0.2825 0.7105 0.3995 0.767 ;
              RECT  0.3425 0.5265 0.3995 0.767 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8955 0.5335 3.118 0.629 ;
              RECT  2.9945 0.4415 3.118 0.629 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END DFFRHQX1

MACRO AOI211XL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6925 0.806 0.9155 ;
              RECT  0.7635 0.2015 0.806 0.9155 ;
              RECT  0.4205 0.318 0.806 0.3605 ;
              RECT  0.7105 0.2015 0.806 0.3605 ;
              RECT  0.4205 0.2015 0.463 0.3605 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.3605 0.113 0.7 ;
              RECT  0.042 0.3605 0.113 0.516 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.325 0.4985 ;
              RECT  0.1835 0.431 0.24 0.7 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3955 0.431 0.537 0.4875 ;
              RECT  0.4665 0.431 0.523 0.7 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.431 0.6645 0.7845 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END AOI211XL

MACRO DFFRX2
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.0825 0.647 3.21 0.7845 ;
              RECT  3.0475 0.3995 3.1465 0.4415 ;
              RECT  3.0825 0.647 3.125 0.9225 ;
              RECT  3.0475 0.3995 3.09 0.689 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.729 0.654 2.786 0.7845 ;
              RECT  2.729 0.378 2.7715 0.9225 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.386 0.7105 2.6585 0.767 ;
              RECT  2.443 0.629 2.4995 0.767 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9085 0.6045 1.1985 0.661 ;
              RECT  0.873 0.576 0.965 0.6325 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.7105 0.3145 0.8375 ;
              RECT  0.258 0.576 0.3145 0.8375 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END DFFRX2

MACRO AND4X6
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.312 0.636 2.3545 0.9685 ;
              RECT  1.732 0.636 2.3545 0.6785 ;
              RECT  1.587 0.371 2.2095 0.4135 ;
              RECT  2.167 0.194 2.2095 0.4135 ;
              RECT  2.022 0.5585 2.0785 0.9685 ;
              RECT  2.022 0.371 2.0645 0.9685 ;
              RECT  1.877 0.194 1.9195 0.4135 ;
              RECT  1.732 0.636 1.7745 0.9685 ;
              RECT  1.587 0.194 1.6295 0.4135 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.5795 1.3715 0.7845 ;
              RECT  0.279 0.795 1.3575 0.8375 ;
              RECT  1.315 0.5795 1.3575 0.8375 ;
              RECT  0.279 0.5795 0.3215 0.8375 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.682 1.2445 0.7245 ;
              RECT  1.202 0.5975 1.2445 0.7245 ;
              RECT  0.4665 0.5585 0.523 0.7245 ;
              RECT  0.392 0.59 0.523 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0145 0.4415 1.1065 0.4985 ;
              RECT  0.5935 0.569 1.071 0.6115 ;
              RECT  1.0285 0.4415 1.071 0.6115 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.4275 0.8235 0.484 ;
              RECT  0.608 0.2895 0.6645 0.484 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END AND4X6

MACRO OR2X4
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.424 1.0885 0.516 ;
              RECT  1.032 0.2965 1.0745 0.76 ;
              RECT  0.9895 0.7175 1.032 0.993 ;
              RECT  0.9895 0.2545 1.032 0.339 ;
              RECT  0.689 0.6045 1.0745 0.647 ;
              RECT  0.7175 0.2965 1.0745 0.339 ;
              RECT  0.668 0.2825 0.753 0.325 ;
              RECT  0.689 0.6045 0.7315 0.993 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.523 0.523 0.8375 ;
              RECT  0.4275 0.523 0.523 0.608 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.187 0.424 0.2435 0.5975 ;
              RECT  0.042 0.424 0.2435 0.4805 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OR2X4

MACRO NAND4X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2615 0.721 0.806 0.7635 ;
              RECT  0.735 0.5585 0.806 0.7635 ;
              RECT  0.735 0.3815 0.7775 0.7635 ;
              RECT  0.5585 0.721 0.601 0.919 ;
              RECT  0.2615 0.721 0.304 0.919 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.021 0.5935 0.24 0.6505 ;
              RECT  0.1625 0.4595 0.24 0.6505 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.325 0.3955 0.629 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.1555 0.523 0.5865 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.2895 0.6645 0.643 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END NAND4X1

MACRO AOI2BB2X1
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.339 1.3715 0.516 ;
              RECT  1.2725 0.424 1.329 0.6505 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.318 1.0885 0.6715 ;
        END
    END B1
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.6645 0.3955 0.721 ;
              RECT  0.332 0.5865 0.3955 0.721 ;
              RECT  0.1835 0.6645 0.24 0.7845 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.4595 0.3815 0.516 ;
              RECT  0.325 0.3815 0.3815 0.516 ;
              RECT  0.1835 0.4595 0.24 0.5935 ;
        END
    END A1N
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1595 0.205 1.202 0.7495 ;
              RECT  0.993 0.205 1.202 0.247 ;
              RECT  0.993 0.173 1.0885 0.247 ;
              RECT  1.032 0.1555 1.0885 0.247 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END AOI2BB2X1

MACRO NAND2BXL
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.028 0.509 0.095 0.5655 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.509 0.636 0.5655 0.774 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1445 0.6115 0.219 0.668 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END NAND2BXL

MACRO DFFSX4
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.719 0.424 4.094 0.4665 ;
              RECT  4.0515 0.3815 4.094 0.4665 ;
              RECT  4.009 0.6645 4.0515 0.94 ;
              RECT  3.719 0.6645 4.0515 0.707 ;
              RECT  3.719 0.424 3.7755 0.707 ;
              RECT  3.719 0.3815 3.7615 0.94 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.429 0.6645 3.4715 0.94 ;
              RECT  3.0545 0.3995 3.429 0.4415 ;
              RECT  3.387 0.357 3.429 0.4415 ;
              RECT  3.1395 0.6645 3.4715 0.707 ;
              RECT  3.1535 0.5585 3.21 0.707 ;
              RECT  3.1535 0.3995 3.196 0.707 ;
              RECT  3.1395 0.6645 3.1815 0.94 ;
              RECT  3.0545 0.357 3.097 0.4415 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.485 0.601 2.5275 0.6855 ;
              RECT  2.1635 0.601 2.5275 0.643 ;
              RECT  2.1635 0.5585 2.22 0.6505 ;
              RECT  2.1775 0.2365 2.22 0.6505 ;
              RECT  1.598 0.2365 2.22 0.279 ;
              RECT  1.3715 0.2685 1.64 0.311 ;
              RECT  1.2865 0.265 1.414 0.3075 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.548 0.463 0.6325 ;
              RECT  0.4065 0.431 0.463 0.6325 ;
              RECT  0.325 0.548 0.3815 0.7035 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.431 0.2545 0.7705 ;
              RECT  0.1835 0.431 0.2545 0.6785 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END DFFSX4

MACRO OR3X6
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.424 1.9125 0.4665 ;
              RECT  1.87 0.247 1.9125 0.4665 ;
              RECT  1.757 0.647 1.7995 0.9685 ;
              RECT  1.177 0.647 1.7995 0.689 ;
              RECT  1.598 0.4205 1.6545 0.516 ;
              RECT  1.598 0.4205 1.64 0.689 ;
              RECT  1.58 0.247 1.6225 0.463 ;
              RECT  1.248 0.4205 1.6545 0.463 ;
              RECT  1.467 0.647 1.5095 0.9685 ;
              RECT  1.248 0.247 1.29 0.463 ;
              RECT  1.177 0.647 1.2195 0.9685 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.601 0.6785 0.6575 ;
              RECT  0.4665 0.601 0.523 0.799 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.4875 0.866 0.5725 ;
              RECT  0.7495 0.4875 0.806 0.6505 ;
              RECT  0.3955 0.4875 0.866 0.53 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.94 0.3745 0.9825 0.523 ;
              RECT  0.1835 0.3745 0.9825 0.417 ;
              RECT  0.1835 0.3745 0.24 0.516 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END OR3X6

MACRO AND3X2
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.424 0.9475 0.516 ;
              RECT  0.8905 0.424 0.933 1.004 ;
              RECT  0.8095 0.424 0.9475 0.4665 ;
              RECT  0.8095 0.339 0.852 0.4665 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.59 0.7105 0.682 0.767 ;
              RECT  0.59 0.7105 0.647 1.0285 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.35 0.3955 0.4065 0.5195 ;
              RECT  0.1835 0.3955 0.4065 0.4525 ;
              RECT  0.1835 0.3955 0.24 0.516 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.113 0.735 ;
              RECT  0.0565 0.3955 0.113 0.735 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END AND3X2

MACRO ADDHXL
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.916 0.371 1.9585 0.735 ;
              RECT  1.8805 0.6925 1.937 0.8025 ;
              RECT  1.8805 0.3285 1.923 0.4135 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3075 0.24 0.8695 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5585 0.6115 0.643 ;
              RECT  0.555 0.537 0.6115 0.643 ;
              RECT  0.4665 0.5585 0.523 0.8025 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1345 0.2155 1.2195 0.258 ;
              RECT  0.9085 0.4665 1.177 0.509 ;
              RECT  1.1345 0.2155 1.177 0.509 ;
              RECT  0.9085 0.2155 0.951 0.509 ;
              RECT  0.4665 0.2155 0.951 0.258 ;
              RECT  0.325 0.424 0.509 0.4665 ;
              RECT  0.4665 0.2155 0.509 0.4665 ;
              RECT  0.325 0.424 0.3955 0.516 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END ADDHXL

MACRO DFFRHQX4
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.333 0.5585 2.6445 0.601 ;
              RECT  2.602 0.516 2.6445 0.601 ;
              RECT  2.333 0.2155 2.3755 0.601 ;
              RECT  1.665 0.2155 2.3755 0.258 ;
              RECT  1.3715 0.35 1.7075 0.392 ;
              RECT  1.665 0.2155 1.7075 0.392 ;
              RECT  1.4385 0.35 1.481 0.5055 ;
              RECT  1.3715 0.2155 1.414 0.392 ;
              RECT  1.0465 0.2155 1.414 0.258 ;
              RECT  1.0355 0.2895 1.0885 0.5125 ;
              RECT  1.0465 0.2155 1.0885 0.5125 ;
              RECT  1.032 0.2895 1.0885 0.3815 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.484 0.3955 0.6325 ;
              RECT  0.134 0.484 0.3955 0.5405 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5775 0.4415 3.765 0.6255 ;
              RECT  3.5775 0.403 3.6345 0.6255 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.774 0.346 0.841 0.7105 ;
              RECT  0.4665 0.668 0.841 0.7105 ;
              RECT  0.4665 0.5585 0.523 0.7105 ;
              RECT  0.424 0.7035 0.509 0.7455 ;
              RECT  0.4665 0.346 0.509 0.7455 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END DFFRHQX4

MACRO NAND3XL
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.6925 0.6645 0.866 ;
              RECT  0.615 0.3815 0.6645 0.866 ;
              RECT  0.286 0.781 0.6645 0.8235 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.537 0.5335 0.622 ;
              RECT  0.4665 0.279 0.523 0.622 ;
        END
    END C
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.021 0.5585 0.24 0.7105 ;
              RECT  0.021 0.5195 0.0775 0.7105 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.339 0.3955 0.629 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END NAND3XL

MACRO SEDFFX4
    CLASS CORE ;
    SIZE 5.6565 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.3875 0.3995 4.7195 0.4415 ;
              RECT  4.6775 0.3425 4.7195 0.4415 ;
              RECT  4.6065 0.721 4.6915 0.7635 ;
              RECT  4.426 0.7105 4.649 0.753 ;
              RECT  4.274 0.742 4.483 0.7845 ;
              RECT  4.426 0.6925 4.483 0.7845 ;
              RECT  4.426 0.3995 4.4685 0.7845 ;
              RECT  4.3875 0.3425 4.43 0.4415 ;
        END
    END QN
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.1545 0.5125 5.473 0.555 ;
              RECT  5.275 0.424 5.3315 0.555 ;
              RECT  4.9815 0.562 5.197 0.6045 ;
              RECT  5.1545 0.5125 5.197 0.6045 ;
              RECT  4.9815 0.562 5.0235 0.675 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.2675 0.6255 5.5115 0.767 ;
              RECT  5.2605 0.6925 5.3315 0.7845 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.122 0.5125 4.2 0.654 ;
              RECT  4.122 0.5125 4.179 0.8445 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.3125 0.3605 3.369 0.6785 ;
              RECT  3.277 0.3605 3.369 0.417 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.136 0.4875 3.235 0.6925 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.647 0.5265 0.951 ;
              RECT  0.484 0.3815 0.5265 0.4665 ;
              RECT  0.4525 0.424 0.4945 0.689 ;
              RECT  0.1835 0.4735 0.4945 0.516 ;
              RECT  0.1835 0.424 0.24 0.516 ;
              RECT  0.1835 0.3815 0.2365 0.951 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.6565 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.6565 0.042 ;
        END
    END VSS
END SEDFFX4

MACRO AND4X4
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2335 0.424 1.3715 0.516 ;
              RECT  1.202 0.7705 1.276 1.0465 ;
              RECT  1.2335 0.339 1.276 1.0465 ;
              RECT  0.88 0.3535 1.276 0.3955 ;
              RECT  1.1415 0.339 1.276 0.3955 ;
              RECT  0.912 0.7705 1.276 0.813 ;
              RECT  0.912 0.7705 0.9545 1.0465 ;
              RECT  0.8305 0.339 0.9155 0.3815 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6925 0.806 0.8905 ;
              RECT  0.707 0.5795 0.7635 0.7495 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.3535 0.523 0.707 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.3675 0.3955 0.707 ;
              RECT  0.325 0.3675 0.3955 0.523 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.3605 0.2545 0.516 ;
              RECT  0.1835 0.424 0.24 0.7 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END AND4X4

MACRO OR4X8
    CLASS CORE ;
    SIZE 2.5455 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.326 0.339 2.411 0.3815 ;
              RECT  1.5095 0.35 2.358 0.392 ;
              RECT  2.3015 0.576 2.344 0.951 ;
              RECT  1.4315 0.576 2.344 0.6185 ;
              RECT  2.1635 0.35 2.22 0.6185 ;
              RECT  2.0575 0.3075 2.1 0.392 ;
              RECT  2.0115 0.576 2.054 0.951 ;
              RECT  1.7465 0.339 1.831 0.392 ;
              RECT  1.7215 0.576 1.764 0.951 ;
              RECT  1.4565 0.339 1.541 0.3815 ;
              RECT  1.4315 0.576 1.474 0.951 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.576 1.248 0.6325 ;
              RECT  1.156 0.548 1.23 0.6325 ;
              RECT  0.1905 0.827 1.1985 0.8695 ;
              RECT  1.156 0.548 1.1985 0.8695 ;
              RECT  0.1905 0.6115 0.233 0.8695 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.714 1.085 0.7565 ;
              RECT  1.0425 0.636 1.085 0.7565 ;
              RECT  0.325 0.6505 0.41 0.7565 ;
              RECT  0.325 0.5585 0.3815 0.7565 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4805 0.601 0.965 0.643 ;
              RECT  0.9225 0.4415 0.965 0.643 ;
              RECT  0.873 0.4415 0.965 0.4985 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4805 0.4735 0.8025 0.53 ;
              RECT  0.4805 0.4415 0.682 0.53 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.5455 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.5455 0.042 ;
        END
    END VSS
END OR4X8

MACRO DFFSHQX1
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1695 0.3815 0.212 0.912 ;
              RECT  0.042 0.424 0.212 0.4665 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.277 0.7105 3.369 0.767 ;
              RECT  3.277 0.569 3.334 0.767 ;
              RECT  3.157 0.569 3.334 0.6255 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9875 0.562 3.0865 0.767 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.9655 0.4805 2.008 0.5655 ;
              RECT  1.81 0.4805 2.008 0.523 ;
              RECT  1.81 0.2545 1.8525 0.523 ;
              RECT  0.8905 0.2545 1.8525 0.2965 ;
              RECT  0.8905 0.424 0.9475 0.516 ;
              RECT  0.682 0.643 0.933 0.6855 ;
              RECT  0.8905 0.2545 0.933 0.6855 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END DFFSHQX1

MACRO SDFFSHQX1
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5585 0.523 0.6505 ;
              RECT  0.339 0.5585 0.523 0.615 ;
              RECT  0.339 0.403 0.424 0.4595 ;
              RECT  0.339 0.403 0.3955 0.721 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.285 0.431 4.3555 0.516 ;
              RECT  4.285 0.424 4.3415 0.516 ;
              RECT  3.712 0.449 4.3555 0.5055 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1185 0.576 4.175 0.7245 ;
              RECT  3.9135 0.576 4.175 0.661 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.224 0.4415 3.415 0.548 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1005 0.6185 3.415 0.675 ;
              RECT  3.1005 0.6185 3.295 0.714 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.686 0.647 1.771 0.689 ;
              RECT  1.407 0.7915 1.7285 0.834 ;
              RECT  1.686 0.647 1.7285 0.834 ;
              RECT  1.407 0.7915 1.4495 0.905 ;
              RECT  1.064 0.8625 1.4495 0.905 ;
              RECT  0.7635 0.873 1.1065 0.9155 ;
              RECT  0.7635 0.6185 0.806 0.9155 ;
              RECT  0.7495 0.6925 0.806 0.7845 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END SDFFSHQX1

MACRO SDFFSHQX4
    CLASS CORE ;
    SIZE 5.091 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.8505 0.456 4.9355 0.4985 ;
              RECT  4.8505 0.424 4.907 0.516 ;
              RECT  4.26 0.463 4.907 0.5055 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.465 0.576 4.78 0.6325 ;
              RECT  4.465 0.576 4.5215 0.6715 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.864 0.4415 3.9205 0.6325 ;
              RECT  3.7015 0.4415 3.9205 0.4985 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.56 0.576 3.751 0.6325 ;
              RECT  3.56 0.4275 3.6305 0.6325 ;
              RECT  3.546 0.4275 3.6305 0.484 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1245 0.707 2.2095 0.7495 ;
              RECT  2.1245 0.707 2.167 0.894 ;
              RECT  1.3715 0.852 2.167 0.894 ;
              RECT  1.0465 0.88 1.414 0.9225 ;
              RECT  1.0465 0.59 1.1805 0.6325 ;
              RECT  1.032 0.827 1.0885 0.919 ;
              RECT  1.0465 0.59 1.0885 0.9225 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5975 0.643 0.6395 0.958 ;
              RECT  0.5975 0.3815 0.6395 0.4665 ;
              RECT  0.5655 0.424 0.608 0.6855 ;
              RECT  0.3075 0.456 0.608 0.4985 ;
              RECT  0.3075 0.424 0.3815 0.516 ;
              RECT  0.3075 0.3815 0.35 0.958 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.091 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.091 0.042 ;
        END
    END VSS
END SDFFSHQX4

MACRO TLATNTSCAX2
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.2895 2.3755 0.3745 ;
              RECT  2.305 0.2895 2.3615 0.912 ;
        END
    END ECK
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.318 0.523 0.6715 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.318 0.3815 0.6715 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0705 0.3605 0.141 0.6715 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END TLATNTSCAX2

MACRO XNOR2X4
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.951 0.5265 1.0355 ;
              RECT  0.484 0.233 0.5265 0.318 ;
              RECT  0.4525 0.76 0.4945 0.993 ;
              RECT  0.1835 0.3885 0.4945 0.431 ;
              RECT  0.4525 0.2755 0.4945 0.431 ;
              RECT  0.1835 0.76 0.4945 0.8025 ;
              RECT  0.173 0.3535 0.258 0.3955 ;
              RECT  0.1835 0.6925 0.24 0.8025 ;
              RECT  0.1835 0.6925 0.2365 1.0355 ;
              RECT  0.1835 0.3535 0.226 1.0355 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.428 0.4415 1.4705 0.5265 ;
              RECT  1.2975 0.4415 1.4705 0.4985 ;
              RECT  1.0075 0.5405 1.3185 0.583 ;
              RECT  1.2125 0.5405 1.2975 0.643 ;
              RECT  1.276 0.456 1.3185 0.583 ;
              RECT  1.0075 0.4595 1.05 0.583 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6785 0.502 0.8235 0.767 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END XNOR2X4

MACRO DFFSX2
    CLASS CORE ;
    SIZE 4.2425 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.698 0.403 3.783 0.4595 ;
              RECT  3.719 0.403 3.7755 0.912 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.295 0.3885 3.3515 0.912 ;
              RECT  3.2665 0.3885 3.3515 0.445 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4465 0.53 2.503 0.8835 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.24 0.7845 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.2425 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.2425 0.042 ;
        END
    END VSS
END DFFSX2

MACRO DFFX2
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.715 0.3745 2.7575 0.912 ;
              RECT  2.588 0.456 2.7575 0.4985 ;
              RECT  2.588 0.424 2.6445 0.516 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.3745 2.3615 0.912 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.022 0.3745 2.0785 0.728 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2015 0.661 0.318 0.7175 ;
              RECT  0.2615 0.6325 0.318 0.7175 ;
              RECT  0.166 0.8445 0.258 0.9015 ;
              RECT  0.2015 0.661 0.258 0.9015 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END DFFX2

MACRO SEDFFX2
    CLASS CORE ;
    SIZE 5.515 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.285 0.6925 4.3695 0.7845 ;
              RECT  4.313 0.2825 4.3695 0.7845 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.3815 0.24 0.912 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.25 0.4415 5.349 0.4985 ;
              RECT  4.7195 0.4135 5.2925 0.456 ;
              RECT  4.7195 0.4135 4.8045 0.4595 ;
              RECT  4.7195 0.4135 4.762 0.767 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.8755 0.5265 5.1795 0.583 ;
              RECT  4.8755 0.5265 5.066 0.6325 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.9845 0.431 4.076 0.6925 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.0295 0.576 3.0865 0.894 ;
              RECT  2.9945 0.576 3.0865 0.6325 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.867 0.5935 2.9235 0.7495 ;
              RECT  2.729 0.5935 2.9235 0.6505 ;
              RECT  2.729 0.5335 2.786 0.6505 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.515 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.515 0.042 ;
        END
    END VSS
END SEDFFX2

MACRO ADDFHXL
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN S
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8885 0.424 3.0685 0.516 ;
              RECT  2.8885 0.3605 2.9305 0.993 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2435 0.6505 0.286 0.8555 ;
              RECT  0.042 0.424 0.286 0.4665 ;
              RECT  0.2435 0.3285 0.286 0.4665 ;
              RECT  0.0565 0.6505 0.286 0.6925 ;
              RECT  0.0565 0.424 0.0985 0.6925 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.895 0.682 2.4995 0.7245 ;
              RECT  1.2055 0.7245 1.937 0.767 ;
              RECT  0.7565 0.682 1.248 0.7245 ;
              RECT  1.149 0.7245 1.937 0.7385 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.57 0.569 2.662 0.6325 ;
              RECT  1.7815 0.569 2.662 0.6115 ;
              RECT  1.3185 0.6115 1.824 0.654 ;
              RECT  0.6395 0.583 1.4035 0.6115 ;
              RECT  0.6395 0.569 1.354 0.6115 ;
              RECT  0.6395 0.569 0.682 0.654 ;
        END
    END A
    PIN CI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0815 0.456 2.287 0.4985 ;
              RECT  1.4915 0.456 1.534 0.5405 ;
              RECT  1.0815 0.4415 1.248 0.4985 ;
        END
    END CI
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END ADDFHXL

MACRO OAI221X2
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.725 0.5585 1.796 0.6505 ;
              RECT  0.4665 0.8165 1.7675 0.859 ;
              RECT  1.725 0.3355 1.7675 0.859 ;
              RECT  1.6545 0.8165 1.697 0.993 ;
              RECT  1.1875 0.8165 1.23 0.9015 ;
              RECT  0.4665 0.8165 0.509 0.9015 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.7035 0.707 0.7455 ;
              RECT  0.6645 0.5975 0.707 0.7455 ;
              RECT  0.1975 0.5585 0.24 0.7455 ;
              RECT  0.1555 0.608 0.24 0.6505 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9895 0.7035 1.513 0.7455 ;
              RECT  1.4565 0.5585 1.513 0.7455 ;
              RECT  0.9895 0.5975 1.032 0.7455 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.449 0.576 0.5935 0.6325 ;
              RECT  0.449 0.5055 0.5055 0.6325 ;
              RECT  0.311 0.5055 0.5055 0.562 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.191 0.5055 1.3855 0.562 ;
              RECT  1.103 0.576 1.248 0.6325 ;
              RECT  1.191 0.5055 1.248 0.6325 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.392 1.6545 0.7455 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END OAI221X2

MACRO SEDFFHQX2
    CLASS CORE ;
    SIZE 4.808 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.668 2.3085 0.7245 ;
              RECT  2.1635 0.35 2.252 0.4065 ;
              RECT  2.1635 0.35 2.22 0.7245 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.582 0.5585 4.787 0.6785 ;
              RECT  4.582 0.4735 4.6385 0.6785 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.036 0.4985 2.093 0.8375 ;
              RECT  2.022 0.4985 2.093 0.6505 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.149 0.4415 1.255 0.6325 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.4135 0.523 0.767 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.636 0.3005 0.6785 0.463 ;
              RECT  0.3535 0.3005 0.6785 0.3425 ;
              RECT  0.166 0.4415 0.3955 0.484 ;
              RECT  0.3535 0.3005 0.3955 0.484 ;
              RECT  0.166 0.4415 0.258 0.4985 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.808 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.808 0.042 ;
        END
    END VSS
END SEDFFHQX2

MACRO SDFFTRX1
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6645 0.2895 0.707 0.94 ;
              RECT  0.608 0.2895 0.707 0.3815 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.912 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.147 0.424 4.3415 0.5195 ;
              RECT  4.285 0.304 4.3415 0.5195 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.9735 0.576 4.076 0.6325 ;
              RECT  3.9735 0.325 4.0305 0.6325 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.6695 0.4415 3.903 0.4985 ;
              RECT  3.6695 0.4415 3.7935 0.6185 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.729 0.555 2.9305 0.6505 ;
              RECT  2.729 0.4415 2.786 0.6505 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7775 0.7105 0.965 0.767 ;
              RECT  0.9085 0.544 0.965 0.767 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END SDFFTRX1

MACRO AND4X2
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9895 0.424 1.0885 0.516 ;
              RECT  0.9225 0.576 1.032 0.6185 ;
              RECT  0.9895 0.251 1.032 0.6185 ;
              RECT  0.9225 0.251 1.032 0.293 ;
              RECT  0.9225 0.576 0.965 0.9435 ;
              RECT  0.9225 0.2085 0.965 0.293 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.548 0.806 0.788 ;
              RECT  0.707 0.477 0.7635 0.6505 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.424 0.523 0.7775 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0245 0.4415 0.2545 0.7035 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END AND4X2

MACRO OAI22XL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.449 0.318 0.562 0.3605 ;
              RECT  0.5195 0.2755 0.562 0.3605 ;
              RECT  0.339 0.4525 0.491 0.4945 ;
              RECT  0.449 0.318 0.491 0.4945 ;
              RECT  0.339 0.4525 0.3815 0.873 ;
              RECT  0.325 0.6925 0.3815 0.7845 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.205 0.41 0.2615 0.6505 ;
              RECT  0.1835 0.5585 0.24 0.742 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.424 0.0985 0.7775 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.431 0.6645 0.7845 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5655 0.523 0.919 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OAI22XL

MACRO DFFSHQX4
    CLASS CORE ;
    SIZE 3.9595 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.7015 0.576 3.7935 0.6325 ;
              RECT  3.737 0.3145 3.7935 0.6325 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1005 0.576 3.3835 0.6325 ;
              RECT  3.1005 0.5055 3.157 0.6325 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1315 0.364 2.174 0.4945 ;
              RECT  1.9445 0.364 2.174 0.4065 ;
              RECT  1.9445 0.251 1.9865 0.4065 ;
              RECT  1.315 0.251 1.9865 0.293 ;
              RECT  1.315 0.424 1.3715 0.516 ;
              RECT  1.0215 0.6115 1.3575 0.654 ;
              RECT  1.315 0.251 1.3575 0.654 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5055 0.3815 0.548 1.0355 ;
              RECT  0.1835 0.4735 0.548 0.516 ;
              RECT  0.2155 0.3815 0.258 1.0355 ;
              RECT  0.1835 0.424 0.258 0.516 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.9595 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.9595 0.042 ;
        END
    END VSS
END DFFSHQX4

MACRO NOR2XL
    CLASS CORE ;
    SIZE 0.5655 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.403 0.8095 ;
              RECT  0.3605 0.304 0.403 0.8095 ;
              RECT  0.1835 0.304 0.403 0.346 ;
              RECT  0.1835 0.2615 0.226 0.346 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.2895 0.113 0.629 ;
              RECT  0.042 0.2895 0.113 0.3815 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.233 0.417 0.2895 0.615 ;
              RECT  0.1835 0.5585 0.24 0.721 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.424 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.424 0.042 ;
        END
    END VSS
END NOR2XL

MACRO XNOR2X2
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2965 0.735 0.3815 0.7915 ;
              RECT  0.325 0.3815 0.3815 0.7915 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.124 0.576 1.4775 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4525 0.576 0.714 0.6325 ;
              RECT  0.4525 0.484 0.6395 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END XNOR2X2

MACRO INVX1
    CLASS CORE ;
    SIZE 0.2825 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.18 0.509 0.2365 0.5655 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0385 0.509 0.1095 0.5655 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.2825 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.2825 0.042 ;
        END
    END VSS
END INVX1

MACRO NAND2X8
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2085 0.742 2.22 0.7845 ;
              RECT  2.1775 0.385 2.22 0.7845 ;
              RECT  2.1635 0.6925 2.22 0.7845 ;
              RECT  0.332 0.385 2.22 0.4275 ;
              RECT  1.948 0.742 1.9905 1.018 ;
              RECT  1.658 0.742 1.7005 1.018 ;
              RECT  1.368 0.742 1.4105 1.018 ;
              RECT  1.078 0.742 1.1205 1.018 ;
              RECT  0.788 0.742 0.8305 1.018 ;
              RECT  0.4985 0.742 0.5405 1.018 ;
              RECT  0.2085 0.7035 0.251 1.018 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.863 0.576 2.0325 0.6185 ;
              RECT  0.53 0.629 1.955 0.6715 ;
              RECT  1.863 0.576 1.955 0.6715 ;
              RECT  1.446 0.6115 1.5305 0.6715 ;
              RECT  1.011 0.6115 1.096 0.6715 ;
              RECT  0.378 0.6115 0.5725 0.654 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.6015 0.516 1.7745 0.5585 ;
              RECT  0.166 0.4985 1.644 0.5405 ;
              RECT  1.255 0.4985 1.3395 0.5585 ;
              RECT  0.643 0.4985 0.728 0.5585 ;
              RECT  0.166 0.4415 0.258 0.5585 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END NAND2X8

MACRO SDFFQX4
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1925 0.456 3.652 0.4985 ;
              RECT  3.56 0.4415 3.652 0.4985 ;
              RECT  3.15 0.654 3.235 0.6965 ;
              RECT  3.1925 0.456 3.235 0.6965 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4185 0.569 3.68 0.6325 ;
              RECT  3.4185 0.569 3.493 0.7175 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.8315 0.5335 3.079 0.6185 ;
              RECT  2.8885 0.5335 2.945 0.6965 ;
              RECT  2.8315 0.5335 2.945 0.6325 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3535 0.24 0.516 ;
              RECT  0.1625 0.4595 0.219 0.6855 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6185 0.403 0.7565 0.445 ;
              RECT  0.6505 0.6255 0.6925 0.912 ;
              RECT  0.6185 0.403 0.661 0.668 ;
              RECT  0.325 0.424 0.661 0.4665 ;
              RECT  0.339 0.403 0.424 0.4665 ;
              RECT  0.3605 0.403 0.403 0.912 ;
              RECT  0.325 0.424 0.403 0.516 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END SDFFQX4

MACRO SDFFXL
    CLASS CORE ;
    SIZE 4.101 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.3815 0.788 0.438 ;
              RECT  0.7315 0.3535 0.788 0.438 ;
              RECT  0.608 0.3815 0.6645 0.8555 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.159 0.2895 0.2155 0.721 ;
              RECT  0.042 0.2895 0.2155 0.449 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.394 0.4415 3.8075 0.4985 ;
              RECT  3.765 0.4135 3.8075 0.4985 ;
              RECT  3.394 0.4135 3.6095 0.4985 ;
              RECT  3.394 0.4135 3.4365 0.6325 ;
              RECT  3.3795 0.59 3.422 0.714 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.7015 0.569 3.8075 0.6785 ;
              RECT  3.507 0.569 3.8075 0.6325 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1395 0.555 3.196 0.6785 ;
              RECT  3.012 0.555 3.196 0.6505 ;
              RECT  3.012 0.4805 3.0685 0.6785 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9085 0.622 1.0005 0.6785 ;
              RECT  0.735 0.7105 0.965 0.767 ;
              RECT  0.9085 0.622 0.965 0.767 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.101 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.101 0.042 ;
        END
    END VSS
END SDFFXL

MACRO CLKBUFX20
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3685 0.647 2.411 0.9615 ;
              RECT  0.042 0.4205 2.411 0.463 ;
              RECT  2.3685 0.251 2.411 0.463 ;
              RECT  0.042 0.647 2.411 0.689 ;
              RECT  2.0785 0.647 2.121 0.9615 ;
              RECT  2.0785 0.251 2.121 0.463 ;
              RECT  1.7885 0.647 1.831 0.9615 ;
              RECT  1.7885 0.251 1.831 0.463 ;
              RECT  1.499 0.647 1.541 0.9615 ;
              RECT  1.499 0.251 1.541 0.463 ;
              RECT  1.209 0.647 1.2515 0.9615 ;
              RECT  1.209 0.251 1.2515 0.463 ;
              RECT  0.919 0.647 0.9615 0.9615 ;
              RECT  0.919 0.251 0.9615 0.463 ;
              RECT  0.629 0.647 0.6715 0.9615 ;
              RECT  0.629 0.251 0.6715 0.463 ;
              RECT  0.339 0.647 0.3815 0.9615 ;
              RECT  0.339 0.251 0.3815 0.463 ;
              RECT  0.042 0.4205 0.0985 0.689 ;
              RECT  0.042 0.251 0.0915 0.9615 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.74 0.576 3.0935 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END CLKBUFX20

MACRO OAI2BB2X2
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8915 0.2825 1.9865 0.325 ;
              RECT  1.467 0.41 1.9335 0.4525 ;
              RECT  1.8915 0.2825 1.9335 0.4525 ;
              RECT  1.7465 0.852 1.7885 0.9365 ;
              RECT  1.467 0.852 1.7885 0.894 ;
              RECT  1.612 0.2825 1.697 0.325 ;
              RECT  1.612 0.2825 1.6545 0.4525 ;
              RECT  1.467 0.41 1.5095 0.894 ;
              RECT  1.0145 0.7245 1.5095 0.767 ;
              RECT  1.1595 0.7245 1.202 1.0285 ;
              RECT  1.0145 0.7105 1.1065 0.767 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.863 0.523 2.008 0.668 ;
              RECT  1.743 0.576 2.008 0.6325 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.58 0.7385 2.121 0.781 ;
              RECT  2.0785 0.615 2.121 0.781 ;
              RECT  1.58 0.576 1.672 0.6325 ;
              RECT  1.58 0.548 1.6225 0.781 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.293 0.576 0.5125 0.6325 ;
              RECT  0.456 0.4415 0.5125 0.6325 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.4415 0.385 0.4985 ;
              RECT  0.166 0.4415 0.2225 0.6325 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END OAI2BB2X2

MACRO FILL32
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END FILL32

MACRO OAI33X1
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.555 0.8555 1.0885 0.898 ;
              RECT  1.018 0.6925 1.0885 0.898 ;
              RECT  1.018 0.2615 1.0605 0.898 ;
              RECT  0.7 0.318 1.0605 0.3605 ;
              RECT  0.9895 0.2615 1.0605 0.3605 ;
              RECT  0.7 0.2615 0.742 0.3605 ;
              RECT  0.555 0.8555 0.5975 1.032 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.431 0.3815 0.7845 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.431 0.6645 0.7845 ;
        END
    END B2
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.24 0.7845 ;
        END
    END A0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.431 0.523 0.7845 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.431 0.806 0.7845 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.431 0.9475 0.7845 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END OAI33X1

MACRO SDFFTRX4
    CLASS CORE ;
    SIZE 5.374 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4335 0.3425 4.8505 0.385 ;
              RECT  4.7305 0.636 4.7725 0.912 ;
              RECT  4.426 0.636 4.7725 0.6785 ;
              RECT  4.426 0.5585 4.483 0.912 ;
              RECT  4.4335 0.3425 4.483 0.912 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1505 0.636 4.193 0.912 ;
              RECT  3.7685 0.3425 4.186 0.385 ;
              RECT  3.8605 0.636 4.193 0.6785 ;
              RECT  3.8745 0.3425 3.917 0.6785 ;
              RECT  3.8605 0.5585 3.903 0.912 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.5585 1.6545 0.7105 ;
              RECT  1.5835 0.371 1.64 0.615 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4565 0.5585 1.513 0.6785 ;
              RECT  1.4105 0.371 1.467 0.615 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.615 0.576 0.8235 0.643 ;
              RECT  0.668 0.4415 0.8235 0.643 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4875 0.4415 0.544 0.7565 ;
              RECT  0.449 0.4415 0.544 0.5265 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.265 0.615 ;
              RECT  0.2085 0.463 0.265 0.615 ;
              RECT  0.042 0.5585 0.0985 0.6505 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.374 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.374 0.042 ;
        END
    END VSS
END SDFFTRX4

MACRO NOR2BXL
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.339 0.279 0.3815 ;
              RECT  0.2365 0.2015 0.279 0.3815 ;
              RECT  0.1625 0.8765 0.205 0.9615 ;
              RECT  0.042 0.8765 0.205 0.919 ;
              RECT  0.042 0.827 0.0985 0.919 ;
              RECT  0.0565 0.339 0.0985 0.919 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.456 0.7495 ;
              RECT  0.3995 0.5055 0.456 0.7495 ;
              RECT  0.325 0.6925 0.3815 0.7845 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.4525 0.24 0.806 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END NOR2BXL

MACRO MXI2X1
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.3425 0.6045 0.385 ;
              RECT  0.4665 0.5585 0.523 0.6505 ;
              RECT  0.4665 0.3425 0.509 0.965 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.82 0.4415 0.965 0.5055 ;
              RECT  0.5865 0.456 0.965 0.4985 ;
              RECT  0.675 0.2295 0.7175 0.4985 ;
              RECT  0.3535 0.2295 0.7175 0.272 ;
              RECT  0.3535 0.2295 0.3955 0.661 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.707 0.576 0.997 0.6325 ;
              RECT  0.707 0.576 0.806 0.6965 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.378 0.24 0.7315 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END MXI2X1

MACRO NOR4BBX1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6925 0.806 0.7845 ;
              RECT  0.3285 0.951 0.7915 0.993 ;
              RECT  0.7495 0.3005 0.7915 0.993 ;
              RECT  0.47 0.3425 0.7915 0.385 ;
              RECT  0.4205 0.3285 0.5055 0.371 ;
              RECT  0.3285 0.951 0.371 1.0355 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.35 0.569 0.424 0.654 ;
              RECT  0.325 0.5975 0.3815 0.88 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.6925 0.6645 0.8095 ;
              RECT  0.4945 0.6925 0.6645 0.7495 ;
              RECT  0.4945 0.569 0.5515 0.7495 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.576 1.1065 0.7565 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0565 0.325 0.113 0.629 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END BN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END NOR4BBX1

MACRO CLKINVX2
    CLASS CORE ;
    SIZE 0.5655 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.3675 0.3815 0.912 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1975 0.424 0.2545 0.5655 ;
              RECT  0.042 0.4805 0.2545 0.537 ;
              RECT  0.042 0.424 0.0985 0.537 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.5655 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.5655 0.042 ;
        END
    END VSS
END CLKINVX2

MACRO SDFFQX2
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2155 0.2615 0.258 0.912 ;
              RECT  0.1835 0.424 0.258 0.516 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.669 0.456 3.1675 0.4985 ;
              RECT  2.853 0.4415 2.945 0.4985 ;
              RECT  2.669 0.456 2.7115 0.5975 ;
              RECT  2.6515 0.555 2.694 0.6785 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.136 0.569 3.2595 0.689 ;
              RECT  2.9695 0.569 3.2595 0.6325 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.5585 2.4675 0.6505 ;
              RECT  2.305 0.4415 2.3615 0.689 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.431 0.523 0.7845 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END SDFFQX2

MACRO AOI22X1
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.661 0.742 0.7035 0.841 ;
              RECT  0.4665 0.742 0.7035 0.7845 ;
              RECT  0.4665 0.6925 0.523 0.7845 ;
              RECT  0.4805 0.2615 0.523 0.7845 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.318 0.806 0.6715 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.2895 0.6645 0.643 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.1905 0.3955 0.4945 ;
              RECT  0.325 0.1555 0.3815 0.247 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END AOI22X1

MACRO TLATNTSCAX20
    CLASS CORE ;
    SIZE 6.2225 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  6.0385 0.537 6.081 0.958 ;
              RECT  6.0385 0.251 6.081 0.4665 ;
              RECT  6.0065 0.424 6.049 0.5795 ;
              RECT  3.719 0.537 6.081 0.5795 ;
              RECT  5.7485 0.251 5.791 0.9615 ;
              RECT  5.4585 0.251 5.501 0.9615 ;
              RECT  5.1685 0.251 5.211 0.9615 ;
              RECT  4.879 0.251 4.921 0.9615 ;
              RECT  4.589 0.251 4.6315 0.9615 ;
              RECT  4.299 0.537 4.3415 0.9615 ;
              RECT  4.299 0.251 4.3415 0.4665 ;
              RECT  4.267 0.424 4.3095 0.5795 ;
              RECT  4.009 0.251 4.0515 0.9615 ;
              RECT  3.719 0.537 3.7755 0.9615 ;
              RECT  3.719 0.251 3.7615 0.9615 ;
        END
    END ECK
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.491 0.576 0.742 0.6325 ;
              RECT  0.523 0.4735 0.682 0.6325 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.364 0.3605 0.4205 0.615 ;
              RECT  0.325 0.5585 0.3815 0.675 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0845 0.4945 0.141 0.7495 ;
              RECT  0.042 0.6925 0.0985 0.806 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.2225 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.2225 0.042 ;
        END
    END VSS
END TLATNTSCAX20

MACRO AO21XL
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.643 0.9155 0.7 ;
              RECT  0.7495 0.286 0.806 0.7 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.5585 0.113 0.7635 ;
              RECT  0.0565 0.424 0.113 0.7635 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5585 0.3675 0.615 ;
              RECT  0.311 0.424 0.3675 0.615 ;
              RECT  0.1835 0.5585 0.24 0.6505 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.516 0.523 0.841 ;
              RECT  0.438 0.516 0.523 0.5725 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END AO21XL

MACRO OAI32XL
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.781 0.523 0.919 0.5655 ;
              RECT  0.8765 0.293 0.919 0.5655 ;
              RECT  0.781 0.523 0.8235 0.873 ;
              RECT  0.7315 0.7105 0.8235 0.767 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.431 0.24 0.7845 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.5585 0.3955 0.898 ;
              RECT  0.325 0.5585 0.3955 0.6505 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.894 0.728 1.0885 0.7845 ;
              RECT  1.032 0.661 1.0885 0.7845 ;
              RECT  0.894 0.636 0.951 0.7845 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.523 0.7105 0.5795 ;
              RECT  0.4665 0.523 0.523 0.689 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.509 1.23 0.6505 ;
              RECT  1.0075 0.509 1.23 0.5655 ;
              RECT  1.0075 0.463 1.064 0.5655 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OAI32XL

MACRO NOR3XL
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.357 0.6645 0.516 ;
              RECT  0.608 0.357 0.6505 0.8305 ;
              RECT  0.5935 0.788 0.636 0.873 ;
              RECT  0.286 0.4945 0.6505 0.537 ;
              RECT  0.286 0.357 0.3285 0.537 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.47 0.608 0.5265 0.7175 ;
              RECT  0.4665 0.661 0.523 0.958 ;
        END
    END C
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.021 0.675 0.2545 0.7845 ;
              RECT  0.021 0.608 0.0775 0.7845 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.668 0.3815 1.0215 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END NOR3XL

MACRO EDFFTRXL
    CLASS CORE ;
    SIZE 4.808 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.3675 0.6645 0.721 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1445 0.3815 0.2015 0.721 ;
              RECT  0.042 0.424 0.2015 0.516 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.426 0.5195 4.55 0.7845 ;
              RECT  4.405 0.5195 4.55 0.6045 ;
        END
    END D
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1255 0.5405 4.2175 0.6325 ;
              RECT  3.8215 0.5405 4.2175 0.5975 ;
        END
    END E
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1535 0.601 3.21 0.834 ;
              RECT  3.033 0.601 3.21 0.6575 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.767 0.4875 0.8235 0.721 ;
              RECT  0.7495 0.385 0.806 0.544 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.808 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.808 0.042 ;
        END
    END VSS
END EDFFTRXL

MACRO MX4X2
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1805 0.3005 1.237 0.4805 ;
              RECT  1.131 0.6785 1.23 0.735 ;
              RECT  1.1735 0.424 1.23 0.735 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.295 0.5585 3.3515 0.6505 ;
              RECT  3.295 0.417 3.3375 0.6505 ;
              RECT  2.8565 0.417 3.3375 0.4595 ;
              RECT  2.8565 0.417 2.899 0.502 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9695 0.53 3.224 0.6325 ;
              RECT  2.9695 0.53 3.026 0.6855 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.3475 0.5935 2.404 0.7495 ;
              RECT  2.305 0.6925 2.3615 0.905 ;
        END
    END C
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.022 0.682 2.121 0.905 ;
              RECT  2.0645 0.5935 2.121 0.905 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.5585 1.5375 0.615 ;
              RECT  1.481 0.463 1.5375 0.615 ;
              RECT  1.315 0.5585 1.3715 0.6505 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.325 0.9475 0.516 ;
              RECT  0.827 0.438 0.898 0.615 ;
        END
    END S1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END MX4X2

MACRO NAND2X6
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.743 0.7175 1.9515 0.767 ;
              RECT  1.909 0.35 1.9515 0.767 ;
              RECT  1.8805 0.6925 1.937 0.7845 ;
              RECT  0.4525 0.35 1.9515 0.392 ;
              RECT  1.743 0.7175 1.785 0.951 ;
              RECT  0.286 0.7175 1.9515 0.76 ;
              RECT  1.527 0.3075 1.5695 0.392 ;
              RECT  1.453 0.7175 1.4955 0.951 ;
              RECT  1.163 0.7175 1.2055 0.951 ;
              RECT  1.0885 0.3075 1.131 0.392 ;
              RECT  0.873 0.7175 0.9155 0.951 ;
              RECT  0.576 0.7175 0.6185 0.951 ;
              RECT  0.4525 0.3075 0.4945 0.392 ;
              RECT  0.286 0.7175 0.3285 0.951 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.576 1.545 0.6325 ;
              RECT  0.647 0.6045 1.474 0.647 ;
              RECT  1.0215 0.576 1.1065 0.647 ;
              RECT  0.502 0.576 0.689 0.6185 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.796 0.463 1.838 0.622 ;
              RECT  0.325 0.463 1.838 0.5055 ;
              RECT  1.2405 0.463 1.3255 0.5265 ;
              RECT  0.76 0.463 0.8445 0.5335 ;
              RECT  0.2435 0.491 0.3815 0.5335 ;
              RECT  0.325 0.424 0.3815 0.5335 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END NAND2X6

MACRO AOI21XL
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.424 0.6645 0.516 ;
              RECT  0.608 0.403 0.6505 0.9155 ;
              RECT  0.5935 0.873 0.636 0.958 ;
              RECT  0.4525 0.403 0.6505 0.445 ;
              RECT  0.4525 0.286 0.4945 0.445 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.431 0.2545 0.4875 ;
              RECT  0.042 0.424 0.0985 0.622 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.1555 0.3815 0.509 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.516 0.523 0.8695 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END AOI21XL

MACRO NAND2X4
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.24 0.7035 1.248 0.7455 ;
              RECT  1.2055 0.35 1.248 0.7455 ;
              RECT  1.156 0.576 1.248 0.6325 ;
              RECT  0.4945 0.35 1.248 0.392 ;
              RECT  1.11 0.7035 1.1525 0.951 ;
              RECT  0.8835 0.3355 0.9685 0.392 ;
              RECT  0.82 0.7035 0.8625 0.951 ;
              RECT  0.53 0.7035 0.5725 0.951 ;
              RECT  0.445 0.3355 0.53 0.378 ;
              RECT  0.24 0.7035 0.2825 0.951 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.456 0.576 0.9155 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.463 1.1345 0.5055 ;
              RECT  0.166 0.4415 0.258 0.5055 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END NAND2X4

MACRO NOR4BBX4
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.005 0.6925 3.0475 0.919 ;
              RECT  2.715 0.6925 3.0475 0.735 ;
              RECT  2.715 0.318 3.0015 0.3605 ;
              RECT  2.959 0.2615 3.0015 0.3605 ;
              RECT  2.715 0.6925 2.786 0.7845 ;
              RECT  2.715 0.2965 2.7575 0.919 ;
              RECT  0.887 0.2965 2.7575 0.339 ;
              RECT  2.669 0.2545 2.7115 0.339 ;
              RECT  2.358 0.2545 2.4005 0.339 ;
              RECT  2.068 0.2545 2.1105 0.339 ;
              RECT  1.757 0.2545 1.7995 0.339 ;
              RECT  1.467 0.2545 1.5095 0.339 ;
              RECT  1.177 0.2545 1.2195 0.339 ;
              RECT  0.887 0.2545 0.9295 0.339 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.588 0.431 2.6445 0.7845 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.022 0.41 2.0785 0.7635 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.537 0.3815 0.8905 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.537 0.24 0.8905 ;
        END
    END BN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END NOR4BBX4

MACRO SDFFSRXL
    CLASS CORE ;
    SIZE 5.374 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.661 0.364 0.7035 0.449 ;
              RECT  0.622 0.3885 0.6645 0.887 ;
              RECT  0.608 0.424 0.6645 0.516 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1625 0.636 0.219 0.721 ;
              RECT  0.1625 0.286 0.219 0.438 ;
              RECT  0.127 0.3745 0.1835 0.7 ;
              RECT  0.042 0.424 0.1835 0.516 ;
              RECT  0.113 0.3745 0.1835 0.516 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.748 0.463 5.2075 0.5055 ;
              RECT  5.1155 0.4415 5.2075 0.5055 ;
              RECT  5.144 0.4205 5.1865 0.5055 ;
              RECT  4.8755 0.4205 4.9175 0.5055 ;
              RECT  4.748 0.463 4.7905 0.707 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.974 0.576 5.144 0.6965 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.5075 0.576 4.564 0.8305 ;
              RECT  4.4085 0.576 4.564 0.6325 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.0835 0.7105 4.437 0.767 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.828 0.9475 3.171 0.9895 ;
              RECT  2.828 0.834 2.8705 0.9895 ;
              RECT  2.1845 0.834 2.8705 0.8765 ;
              RECT  2.1845 0.6715 2.227 0.8765 ;
              RECT  1.6295 0.6715 2.227 0.714 ;
              RECT  1.6295 0.576 1.672 0.714 ;
              RECT  1.4845 0.59 1.672 0.6325 ;
              RECT  1.58 0.576 1.672 0.6325 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.88 0.7035 0.9825 0.799 ;
              RECT  0.735 0.636 0.965 0.767 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.374 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.374 0.042 ;
        END
    END VSS
END SDFFSRXL

MACRO OR3X1
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.2615 0.806 0.919 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.449 0.4415 0.5655 0.735 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2085 0.456 0.265 0.7845 ;
              RECT  0.1835 0.456 0.265 0.6505 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.431 0.0985 0.7845 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OR3X1

MACRO AOI211X2
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.156 0.3145 1.2405 0.357 ;
              RECT  1.177 0.668 1.2195 0.866 ;
              RECT  0.438 0.3285 1.191 0.371 ;
              RECT  0.7635 0.668 1.2195 0.7105 ;
              RECT  0.8445 0.3145 0.9295 0.371 ;
              RECT  0.7635 0.3285 0.806 0.7105 ;
              RECT  0.7495 0.3285 0.806 0.516 ;
              RECT  0.3885 0.3145 0.4735 0.357 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.371 0.569 0.6325 0.647 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.4415 0.6395 0.4985 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0145 0.4415 1.131 0.5975 ;
              RECT  0.8765 0.4415 1.131 0.4985 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.202 0.4415 1.389 0.562 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END AOI211X2

MACRO BUFX6
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.403 1.0885 0.7565 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.629 0.647 0.6715 0.9685 ;
              RECT  0.042 0.4205 0.6715 0.463 ;
              RECT  0.629 0.247 0.6715 0.463 ;
              RECT  0.042 0.647 0.6715 0.689 ;
              RECT  0.339 0.647 0.3815 0.9685 ;
              RECT  0.339 0.247 0.3815 0.463 ;
              RECT  0.042 0.5585 0.0985 0.689 ;
              RECT  0.042 0.247 0.0915 0.9685 ;
        END
    END Y
END BUFX6

MACRO NOR3BXL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.357 0.2155 0.4525 0.258 ;
              RECT  0.0565 0.332 0.3995 0.3745 ;
              RECT  0.357 0.2155 0.3995 0.3745 ;
              RECT  0.152 0.8695 0.194 0.9545 ;
              RECT  0.0565 0.8695 0.194 0.912 ;
              RECT  0.0985 0.194 0.141 0.3745 ;
              RECT  0.0565 0.332 0.0985 0.912 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5405 0.548 0.682 0.6325 ;
              RECT  0.583 0.53 0.6395 0.6325 ;
              RECT  0.5405 0.548 0.5975 0.799 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.445 0.3815 0.799 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.445 0.24 0.799 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END NOR3BXL

MACRO MXI3X1
    CLASS CORE ;
    SIZE 2.687 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.588 0.3815 2.6445 0.912 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.438 2.404 0.523 ;
              RECT  2.287 0.438 2.344 0.608 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.58 0.643 1.955 0.7 ;
              RECT  1.58 0.576 1.672 0.7 ;
              RECT  1.58 0.5655 1.665 0.7 ;
        END
    END S1
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.004 0.7105 1.2405 0.767 ;
              RECT  1.004 0.5935 1.0605 0.767 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2615 0.548 0.5795 0.6045 ;
              RECT  0.2615 0.548 0.3995 0.6395 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.134 0.7105 0.707 0.767 ;
              RECT  0.6505 0.6575 0.707 0.767 ;
              RECT  0.134 0.6325 0.1905 0.767 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.687 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.687 0.042 ;
        END
    END VSS
END MXI3X1

MACRO NAND2BX2
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.053 0.3885 0.1095 0.449 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7315 0.548 0.788 0.661 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.053 0.675 0.1095 0.7315 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END NAND2BX2

MACRO AOI32X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.781 0.7105 0.8235 0.9225 ;
              RECT  0.601 0.7105 0.8235 0.767 ;
              RECT  0.601 0.357 0.643 0.767 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.339 0.339 0.3955 0.629 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.873 0.4415 0.965 0.4985 ;
              RECT  0.714 0.544 0.9295 0.601 ;
              RECT  0.873 0.4415 0.9295 0.601 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4735 0.325 0.53 0.636 ;
              RECT  0.4665 0.2895 0.523 0.3815 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0355 0.4595 1.23 0.516 ;
              RECT  1.1735 0.424 1.23 0.516 ;
              RECT  1.0355 0.4595 1.092 0.6395 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.4135 0.24 0.767 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END AOI32X1

MACRO OAI2BB1XL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2895 0.8625 0.332 0.9475 ;
              RECT  0.212 0.8625 0.332 0.905 ;
              RECT  0.212 0.438 0.2545 0.905 ;
              RECT  0.0565 0.212 0.24 0.2545 ;
              RECT  0.1975 0.1695 0.24 0.2545 ;
              RECT  0.0565 0.438 0.2545 0.4805 ;
              RECT  0.0565 0.212 0.0985 0.4805 ;
              RECT  0.042 0.2895 0.0985 0.3815 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.438 0.3815 0.7915 ;
        END
    END B0
    PIN A0N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.438 0.523 0.7915 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.431 0.806 0.7845 ;
        END
    END A1N
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END OAI2BB1XL

MACRO AO22XL
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.643 1.0675 0.7 ;
              RECT  0.8905 0.424 0.9475 0.7 ;
              RECT  0.8835 0.286 0.94 0.4805 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.5585 0.806 0.8695 ;
              RECT  0.707 0.5585 0.806 0.615 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.4205 0.523 0.774 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.1625 0.3815 0.516 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END AO22XL

MACRO NAND2X2
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.615 0.537 0.6715 0.5935 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2545 0.438 0.403 0.509 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0455 0.5655 0.106 0.6925 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END NAND2X2

MACRO NOR4XL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.735 0.6925 0.806 0.7845 ;
              RECT  0.7635 0.3425 0.806 0.7845 ;
              RECT  0.247 0.3425 0.806 0.385 ;
              RECT  0.5585 0.205 0.601 0.385 ;
              RECT  0.247 0.205 0.2895 0.385 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.021 0.576 0.2545 0.6325 ;
              RECT  0.088 0.456 0.2545 0.6325 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.516 0.3815 0.8695 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.456 0.523 0.8095 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.4595 0.6925 0.516 ;
              RECT  0.608 0.4595 0.6645 0.7845 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END NOR4XL

MACRO MX3XL
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.028 0.8695 0.113 0.912 ;
              RECT  0.0705 0.2895 0.113 0.912 ;
              RECT  0.042 0.2895 0.113 0.3815 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4315 0.767 1.796 0.8235 ;
              RECT  1.739 0.6925 1.796 0.8235 ;
              RECT  1.4315 0.5865 1.488 0.8235 ;
              RECT  1.389 0.5585 1.446 0.643 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.559 0.523 1.796 0.5795 ;
              RECT  1.598 0.523 1.6545 0.6965 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0355 0.424 1.092 0.7565 ;
              RECT  1.032 0.4065 1.0885 0.548 ;
        END
    END B
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.887 0.6715 0.9475 0.7565 ;
              RECT  0.8905 0.4065 0.9475 0.7565 ;
        END
    END S1
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5405 0.2895 0.6255 ;
              RECT  0.1835 0.5405 0.24 0.8445 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END MX3XL

MACRO CLKINVX8
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.078 0.403 1.163 0.445 ;
              RECT  1.0995 0.6785 1.1415 0.951 ;
              RECT  0.2615 0.4135 1.11 0.456 ;
              RECT  0.8025 0.6785 1.1415 0.721 ;
              RECT  0.8905 0.4135 0.9475 0.516 ;
              RECT  0.8905 0.4135 0.933 0.721 ;
              RECT  0.8095 0.6785 0.852 0.951 ;
              RECT  0.8095 0.371 0.852 0.456 ;
              RECT  0.2295 0.7035 0.852 0.7455 ;
              RECT  0.4985 0.403 0.583 0.456 ;
              RECT  0.5195 0.7035 0.562 0.951 ;
              RECT  0.2085 0.403 0.293 0.445 ;
              RECT  0.2295 0.7035 0.272 0.951 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.544 0.774 0.601 ;
              RECT  0.3075 0.544 0.3995 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END CLKINVX8

MACRO NAND4BX1
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5515 0.8485 0.5935 1.0465 ;
              RECT  0.042 0.8485 0.5935 0.8905 ;
              RECT  0.2545 0.8485 0.2965 1.0465 ;
              RECT  0.0565 0.311 0.187 0.3535 ;
              RECT  0.1445 0.2685 0.187 0.3535 ;
              RECT  0.042 0.6925 0.0985 0.8905 ;
              RECT  0.0565 0.311 0.0985 0.8905 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.537 0.806 0.8905 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4595 0.5585 0.523 0.6505 ;
              RECT  0.4595 0.304 0.516 0.6505 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.332 0.5655 0.3885 0.7775 ;
              RECT  0.325 0.431 0.3815 0.6505 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.24 0.7775 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END NAND4BX1

MACRO AOI31XL
    CLASS CORE ;
    SIZE 1.131 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.894 0.5585 1.0885 0.6505 ;
              RECT  0.894 0.5195 0.9365 0.8555 ;
              RECT  0.636 0.5195 0.9365 0.562 ;
              RECT  0.636 0.3815 0.6785 0.562 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5585 0.24 0.767 ;
              RECT  0.0385 0.5585 0.24 0.6325 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.767 0.6575 0.8235 0.9755 ;
              RECT  0.7315 0.6575 0.8235 0.767 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.509 0.456 0.5655 0.767 ;
              RECT  0.4665 0.456 0.5655 0.6505 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3285 0.3005 0.385 0.643 ;
              RECT  0.325 0.5585 0.3815 0.6505 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.131 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.131 0.042 ;
        END
    END VSS
END AOI31XL

MACRO DLY1X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.3675 1.23 0.912 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.438 0.3815 0.6645 ;
              RECT  0.1975 0.548 0.3815 0.6325 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END DLY1X1

MACRO OAI21X4
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.644 0.3355 1.739 0.378 ;
              RECT  1.3255 0.371 1.686 0.4135 ;
              RECT  1.605 0.7315 1.6475 0.972 ;
              RECT  1.315 0.7315 1.6475 0.774 ;
              RECT  1.3255 0.3355 1.4495 0.4135 ;
              RECT  1.315 0.7315 1.3715 0.919 ;
              RECT  0.445 0.721 1.368 0.7635 ;
              RECT  1.3255 0.3355 1.368 0.919 ;
              RECT  1.315 0.721 1.3575 0.972 ;
              RECT  0.8835 0.721 0.926 0.972 ;
              RECT  0.445 0.721 0.4875 0.972 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.5865 0.894 0.643 ;
              RECT  0.3075 0.576 0.4805 0.643 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.5585 1.23 0.6505 ;
              RECT  1.1135 0.5585 1.23 0.601 ;
              RECT  1.1135 0.463 1.156 0.601 ;
              RECT  0.212 0.463 1.156 0.5055 ;
              RECT  0.59 0.463 0.675 0.516 ;
              RECT  0.148 0.4665 0.2365 0.509 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.4385 0.576 1.672 0.6325 ;
              RECT  1.4385 0.484 1.4955 0.661 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END OAI21X4

MACRO SDFFRHQX8
    CLASS CORE ;
    SIZE 5.515 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.1935 0.4415 5.349 0.5055 ;
              RECT  4.794 0.456 5.349 0.4985 ;
              RECT  4.794 0.456 4.8365 0.647 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.0415 0.576 5.381 0.6325 ;
              RECT  5.0415 0.576 5.2075 0.647 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.5535 0.4415 4.61 0.6325 ;
              RECT  4.426 0.4415 4.61 0.4985 ;
              RECT  4.426 0.424 4.483 0.516 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.404 0.576 2.584 0.647 ;
              RECT  2.5065 0.417 2.584 0.647 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.6895 0.491 1.7995 0.5335 ;
              RECT  1.6895 0.2435 1.732 0.5335 ;
              RECT  1.347 0.2435 1.732 0.286 ;
              RECT  1.276 0.4985 1.389 0.5405 ;
              RECT  1.347 0.2435 1.389 0.5405 ;
              RECT  1.2975 0.4415 1.389 0.5405 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0075 0.424 1.11 0.4665 ;
              RECT  1.0675 0.3815 1.11 0.4665 ;
              RECT  1.0075 0.424 1.05 0.9545 ;
              RECT  0.1375 0.4735 1.05 0.516 ;
              RECT  0.7775 0.3815 0.82 0.516 ;
              RECT  0.7175 0.4735 0.76 0.9545 ;
              RECT  0.4875 0.3815 0.53 0.516 ;
              RECT  0.4275 0.4735 0.47 0.9545 ;
              RECT  0.1835 0.3815 0.24 0.516 ;
              RECT  0.1375 0.4735 0.18 0.9545 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.515 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.515 0.042 ;
        END
    END VSS
END SDFFRHQX8

MACRO NAND4BBX2
    CLASS CORE ;
    SIZE 2.2625 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.096 0.774 2.068 0.8165 ;
              RECT  2.0255 0.311 2.068 0.8165 ;
              RECT  1.994 0.774 2.036 0.972 ;
              RECT  1.6755 0.774 1.718 0.972 ;
              RECT  1.3855 0.774 1.428 0.972 ;
              RECT  1.096 0.7105 1.248 0.8165 ;
              RECT  1.096 0.7105 1.138 0.972 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8985 0.4595 1.955 0.7035 ;
              RECT  1.8805 0.3675 1.937 0.516 ;
        END
    END D
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.5905 0.5585 1.796 0.7035 ;
              RECT  1.5905 0.4985 1.6475 0.7035 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3995 0.7105 0.562 0.8235 ;
              RECT  0.3995 0.576 0.4595 0.8235 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.272 0.576 0.3285 0.8235 ;
              RECT  0.166 0.576 0.3285 0.6325 ;
        END
    END BN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.2625 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.2625 0.042 ;
        END
    END VSS
END NAND4BBX2

MACRO SDFFSXL
    CLASS CORE ;
    SIZE 4.384 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7635 0.403 0.8485 0.4595 ;
              RECT  0.7635 0.403 0.82 0.7035 ;
              RECT  0.7495 0.647 0.806 0.7845 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.403 0.3815 0.516 ;
              RECT  0.325 0.403 0.3675 0.8625 ;
              RECT  0.2965 0.403 0.3815 0.445 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.836 0.456 4.221 0.4985 ;
              RECT  4.1255 0.4415 4.2175 0.4985 ;
              RECT  3.97 0.4135 4.0125 0.4985 ;
              RECT  3.7615 0.682 3.878 0.7245 ;
              RECT  3.836 0.456 3.878 0.7245 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.069 0.576 4.2035 0.7245 ;
              RECT  4.147 0.569 4.2035 0.7245 ;
              RECT  3.949 0.576 4.2035 0.6325 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.521 0.4135 3.652 0.4985 ;
              RECT  3.521 0.4135 3.5775 0.6925 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.3125 0.622 3.4505 0.6785 ;
              RECT  3.3125 0.4415 3.369 0.6785 ;
              RECT  3.277 0.4415 3.369 0.4985 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.916 0.2895 2.227 0.332 ;
              RECT  2.1845 0.247 2.227 0.332 ;
              RECT  1.916 0.205 1.9585 0.332 ;
              RECT  1.488 0.205 1.9585 0.247 ;
              RECT  1.2125 0.576 1.5305 0.6185 ;
              RECT  1.488 0.205 1.5305 0.6185 ;
              RECT  1.2975 0.576 1.389 0.6325 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.384 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.384 0.042 ;
        END
    END VSS
END SDFFSXL

MACRO MX2X4
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.368 0.742 1.4105 1.0465 ;
              RECT  1.11 0.332 1.4105 0.3745 ;
              RECT  1.368 0.2755 1.4105 0.3745 ;
              RECT  1.078 0.742 1.4105 0.7845 ;
              RECT  1.11 0.6925 1.23 0.7845 ;
              RECT  1.11 0.2965 1.1525 0.7845 ;
              RECT  1.078 0.742 1.1205 1.0465 ;
              RECT  1.057 0.2965 1.1525 0.339 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.873 0.576 1.039 0.6325 ;
              RECT  0.834 0.6715 0.9295 0.781 ;
              RECT  0.873 0.576 0.9295 0.781 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.445 0.3815 0.799 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4525 0.643 0.537 0.6855 ;
              RECT  0.1835 0.8695 0.4945 0.912 ;
              RECT  0.4525 0.643 0.4945 0.912 ;
              RECT  0.1835 0.6925 0.24 0.912 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END MX2X4

MACRO NOR4BXL
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.6965 0.205 0.781 0.247 ;
              RECT  0.0565 0.3215 0.7385 0.364 ;
              RECT  0.6965 0.205 0.7385 0.364 ;
              RECT  0.4275 0.1835 0.47 0.364 ;
              RECT  0.3355 0.721 0.378 0.806 ;
              RECT  0.0565 0.721 0.378 0.7635 ;
              RECT  0.0565 0.3215 0.0985 0.7635 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.894 0.576 1.1065 0.6325 ;
              RECT  0.9755 0.4345 1.032 0.6325 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.5585 0.806 0.6925 ;
              RECT  0.654 0.5585 0.806 0.615 ;
              RECT  0.654 0.4345 0.7105 0.615 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.484 0.491 0.583 0.548 ;
              RECT  0.449 0.7105 0.5405 0.767 ;
              RECT  0.484 0.491 0.5405 0.767 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.516 0.378 0.6505 ;
              RECT  0.3215 0.4345 0.378 0.6505 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END NOR4BXL

MACRO MXI4X1
    CLASS CORE ;
    SIZE 2.9695 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0915 0.3815 0.148 0.9475 ;
              RECT  0.042 0.424 0.148 0.516 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4075 0.576 2.761 0.6325 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4075 0.753 2.6795 0.841 ;
              RECT  2.4075 0.7035 2.5205 0.841 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.983 0.6645 2.0965 0.841 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7005 0.7105 1.9125 0.767 ;
              RECT  1.8275 0.569 1.9125 0.767 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.191 0.636 1.4035 0.707 ;
              RECT  1.191 0.576 1.248 0.707 ;
              RECT  1.124 0.576 1.248 0.6325 ;
        END
    END D
    PIN S1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.011 0.173 1.0535 0.622 ;
              RECT  0.7315 0.173 1.0535 0.2155 ;
              RECT  0.339 0.1905 0.774 0.233 ;
              RECT  0.339 0.1905 0.3815 0.5865 ;
              RECT  0.325 0.2895 0.3815 0.3815 ;
        END
    END S1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.9695 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.9695 0.042 ;
        END
    END VSS
END MXI4X1

MACRO OAI21X2
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.424 0.979 0.4665 ;
              RECT  0.9365 0.3815 0.979 0.4665 ;
              RECT  0.456 0.806 0.919 0.8485 ;
              RECT  0.8765 0.424 0.919 0.8485 ;
              RECT  0.8445 0.806 0.887 1.0465 ;
              RECT  0.7495 0.608 0.919 0.6505 ;
              RECT  0.7495 0.5585 0.806 0.6505 ;
              RECT  0.456 0.806 0.4985 1.0465 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6785 0.4945 0.735 ;
              RECT  0.325 0.6785 0.3815 0.919 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.5515 0.6645 0.6505 ;
              RECT  0.2435 0.5515 0.6645 0.608 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9895 0.5585 1.0885 0.6505 ;
              RECT  0.9895 0.537 1.0465 0.8485 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OAI21X2

MACRO NAND4BX4
    CLASS CORE ;
    SIZE 3.111 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.192 0.357 2.8495 0.3995 ;
              RECT  2.807 0.3005 2.8495 0.3995 ;
              RECT  2.6265 0.7035 2.669 0.958 ;
              RECT  1.032 0.7035 2.669 0.7455 ;
              RECT  2.4995 0.3005 2.542 0.3995 ;
              RECT  2.3365 0.7035 2.379 0.958 ;
              RECT  1.0465 0.463 2.234 0.5055 ;
              RECT  2.192 0.357 2.234 0.5055 ;
              RECT  1.9445 0.7035 1.9865 0.958 ;
              RECT  1.6545 0.7035 1.697 0.958 ;
              RECT  1.3645 0.7035 1.407 0.958 ;
              RECT  1.0745 0.7035 1.117 0.958 ;
              RECT  0.484 0.682 1.0885 0.7245 ;
              RECT  1.032 0.7035 1.117 0.7845 ;
              RECT  1.0465 0.463 1.0885 0.7845 ;
              RECT  0.774 0.682 0.8165 0.958 ;
              RECT  0.484 0.682 0.5265 0.958 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0705 0.4595 0.127 0.7495 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1595 0.576 1.513 0.6325 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.305 0.47 2.39 0.5125 ;
              RECT  1.732 0.59 2.3475 0.6325 ;
              RECT  2.305 0.47 2.3475 0.6325 ;
              RECT  2.146 0.576 2.3475 0.6325 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.5595 0.47 2.7715 0.5265 ;
              RECT  2.432 0.576 2.662 0.6325 ;
              RECT  2.5595 0.47 2.662 0.6325 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.111 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.111 0.042 ;
        END
    END VSS
END NAND4BX4

MACRO TIEHI
    CLASS CORE ;
    SIZE 0.424 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.636 0.0985 0.9895 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.424 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.424 0.042 ;
        END
    END VSS
END TIEHI

MACRO CLKINVX12
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.194 0.636 1.5305 0.6785 ;
              RECT  1.488 0.3285 1.5305 0.6785 ;
              RECT  1.4565 0.636 1.513 0.9685 ;
              RECT  0.233 0.3285 1.5305 0.371 ;
              RECT  1.407 0.1625 1.4495 0.371 ;
              RECT  1.103 0.636 1.1455 0.9685 ;
              RECT  1.103 0.1625 1.1455 0.371 ;
              RECT  0.813 0.636 0.8555 0.9685 ;
              RECT  0.813 0.1625 0.8555 0.371 ;
              RECT  0.523 0.636 0.5655 0.9685 ;
              RECT  0.523 0.1625 0.5655 0.371 ;
              RECT  0.233 0.1625 0.2755 0.371 ;
              RECT  0.194 0.636 0.2365 0.9685 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.265 0.4415 1.4175 0.484 ;
              RECT  0.3075 0.4415 0.3995 0.4985 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END CLKINVX12

MACRO OA21X4
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8485 0.6645 1.3715 0.707 ;
              RECT  1.2405 0.5585 1.3715 0.707 ;
              RECT  1.2405 0.438 1.283 0.707 ;
              RECT  1.209 0.3815 1.2515 0.4805 ;
              RECT  0.919 0.438 1.283 0.4805 ;
              RECT  1.138 0.6645 1.1805 0.9545 ;
              RECT  0.919 0.3815 0.9615 0.4805 ;
              RECT  0.8485 0.6645 0.8905 0.9545 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.445 0.0985 0.799 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3075 0.445 0.4275 0.6325 ;
              RECT  0.205 0.445 0.4275 0.502 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.5585 0.6645 0.6855 ;
              RECT  0.509 0.5585 0.6645 0.615 ;
              RECT  0.509 0.431 0.5655 0.615 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END OA21X4

MACRO AOI221XL
    CLASS CORE ;
    SIZE 1.414 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.2865 0.5585 1.3715 0.6505 ;
              RECT  1.2865 0.4525 1.329 0.8555 ;
              RECT  0.682 0.4525 1.329 0.4945 ;
              RECT  1.2125 0.3355 1.255 0.4945 ;
              RECT  0.682 0.3355 0.7245 0.4945 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4875 0.6185 0.799 0.675 ;
              RECT  0.4875 0.576 0.682 0.675 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8695 0.576 1.0885 0.6325 ;
              RECT  0.88 0.576 0.9365 0.767 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.166 0.59 0.279 0.767 ;
        END
    END A0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0075 0.7105 1.216 0.767 ;
              RECT  1.1595 0.5655 1.216 0.767 ;
        END
    END C0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.332 0.463 0.417 0.5195 ;
              RECT  0.332 0.173 0.3995 0.5195 ;
              RECT  0.3075 0.173 0.3995 0.2295 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.414 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.414 0.042 ;
        END
    END VSS
END AOI221XL

MACRO DLY2X1
    CLASS CORE ;
    SIZE 2.404 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1905 0.788 0.233 0.986 ;
              RECT  0.0565 0.293 0.233 0.3355 ;
              RECT  0.1905 0.251 0.233 0.3355 ;
              RECT  0.0565 0.788 0.233 0.8305 ;
              RECT  0.0565 0.293 0.0985 0.8305 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.424 1.0885 0.516 ;
              RECT  1.018 0.4415 1.0745 0.7635 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.404 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.404 0.042 ;
        END
    END VSS
END DLY2X1

MACRO OAI31X4
    CLASS CORE ;
    SIZE 2.828 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.503 0.3425 2.5985 0.385 ;
              RECT  2.1635 0.378 2.5455 0.4205 ;
              RECT  2.464 0.7175 2.5065 0.993 ;
              RECT  2.1635 0.742 2.5065 0.7845 ;
              RECT  2.1635 0.3425 2.3085 0.4205 ;
              RECT  2.1635 0.6925 2.22 0.7845 ;
              RECT  2.174 0.6925 2.2165 0.993 ;
              RECT  2.1635 0.3425 2.206 0.8375 ;
              RECT  0.647 0.795 2.2165 0.8375 ;
              RECT  1.5305 0.795 1.573 0.993 ;
              RECT  0.647 0.795 0.689 0.993 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4215 0.5655 2.6195 0.6325 ;
              RECT  2.2765 0.5655 2.6195 0.622 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4275 0.682 1.994 0.7245 ;
              RECT  1.9515 0.6045 1.994 0.7245 ;
              RECT  1.0075 0.6255 1.092 0.7245 ;
              RECT  0.4275 0.6185 0.47 0.7245 ;
              RECT  0.166 0.6185 0.47 0.661 ;
              RECT  0.166 0.576 0.258 0.661 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.598 0.4415 1.8135 0.5265 ;
              RECT  1.598 0.424 1.6545 0.5265 ;
              RECT  1.163 0.569 1.64 0.6115 ;
              RECT  1.598 0.424 1.64 0.6115 ;
              RECT  1.163 0.5125 1.2055 0.6115 ;
              RECT  0.894 0.5125 1.2055 0.555 ;
              RECT  0.5405 0.569 0.9365 0.6115 ;
              RECT  0.894 0.5125 0.9365 0.6115 ;
              RECT  0.5405 0.463 0.583 0.6115 ;
              RECT  0.3145 0.463 0.583 0.5055 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.276 0.456 1.4955 0.4985 ;
              RECT  1.276 0.3995 1.3185 0.4985 ;
              RECT  0.781 0.3995 1.3185 0.4415 ;
              RECT  0.654 0.456 0.8235 0.4985 ;
              RECT  0.7315 0.4415 0.8235 0.4985 ;
        END
    END A2
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.828 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.828 0.042 ;
        END
    END VSS
END OAI31X4

MACRO TLATNTSCAX12
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.154 0.6715 4.1965 1.004 ;
              RECT  3.012 0.5585 4.1965 0.601 ;
              RECT  4.154 0.247 4.1965 0.601 ;
              RECT  4.122 0.5585 4.1645 0.714 ;
              RECT  3.864 0.247 3.9065 1.004 ;
              RECT  3.574 0.247 3.6165 1.004 ;
              RECT  3.2845 0.247 3.3265 1.004 ;
              RECT  3.012 0.5585 3.0685 0.6505 ;
              RECT  3.012 0.4275 3.0545 0.6505 ;
              RECT  2.9945 0.615 3.0405 0.654 ;
              RECT  2.9945 0.615 3.037 1.004 ;
              RECT  2.9945 0.247 3.037 0.4665 ;
        END
    END ECK
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.47 0.318 0.5265 0.668 ;
              RECT  0.4665 0.318 0.5265 0.516 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.318 0.3815 0.668 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.339 0.0985 0.6325 ;
        END
    END E
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END TLATNTSCAX12

MACRO NAND3BXL
    CLASS CORE ;
    SIZE 0.707 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.042 0.7105 0.0985 0.767 ;
        END
    END Y
    PIN AN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.5125 0.5405 0.5725 0.6325 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.233 0.325 0.3285 0.364 ;
              RECT  0.233 0.2895 0.2895 0.364 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.127 0.424 0.1905 0.4985 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.707 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.707 0.042 ;
        END
    END VSS
END NAND3BXL

MACRO EDFFX4
    CLASS CORE ;
    SIZE 4.525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.9985 0.742 4.041 1.018 ;
              RECT  3.606 0.403 4.023 0.445 ;
              RECT  3.7085 0.742 4.041 0.7845 ;
              RECT  3.719 0.6925 3.7755 0.7845 ;
              RECT  3.719 0.403 3.7615 0.7845 ;
              RECT  3.7085 0.742 3.751 1.018 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4185 0.742 3.461 1.018 ;
              RECT  3.1285 0.742 3.461 0.7845 ;
              RECT  2.9415 0.403 3.3585 0.445 ;
              RECT  3.1535 0.6925 3.21 0.7845 ;
              RECT  3.1535 0.403 3.196 0.7845 ;
              RECT  3.1285 0.742 3.171 1.018 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.577 0.576 2.9305 0.6325 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.153 0.576 2.2375 0.788 ;
              RECT  2.04 0.576 2.2375 0.6325 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5405 0.24 0.894 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.525 0.042 ;
        END
    END VSS
END EDFFX4

MACRO OAI222X1
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.491 0.841 1.23 0.8835 ;
              RECT  1.1735 0.6925 1.23 0.8835 ;
              RECT  1.1735 0.318 1.216 0.8835 ;
              RECT  1.018 0.318 1.216 0.3605 ;
              RECT  1.057 0.841 1.0995 1.039 ;
              RECT  1.018 0.2615 1.0605 0.3605 ;
              RECT  0.491 0.841 0.5335 1.039 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.5585 0.5865 0.7705 ;
              RECT  0.53 0.4805 0.5865 0.7705 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.4805 0.24 0.834 ;
        END
    END A0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8905 0.417 0.9475 0.7705 ;
        END
    END C0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.6925 0.3815 0.82 ;
              RECT  0.311 0.4805 0.3675 0.7495 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.5585 1.103 0.7705 ;
              RECT  1.0465 0.431 1.103 0.7705 ;
        END
    END C1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.318 0.806 0.6715 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OAI222X1

MACRO SDFFRHQX2
    CLASS CORE ;
    SIZE 4.101 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.654 0.24 0.9295 ;
              RECT  0.18 0.2965 0.2365 0.7105 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.6345 0.463 3.871 0.5055 ;
              RECT  3.3795 0.456 3.6765 0.4985 ;
              RECT  3.56 0.4415 3.652 0.4985 ;
              RECT  3.3795 0.456 3.422 0.647 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.6345 0.5975 3.9665 0.654 ;
              RECT  3.673 0.576 3.9665 0.654 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.1395 0.424 3.196 0.615 ;
              RECT  3.012 0.424 3.196 0.4805 ;
              RECT  3.012 0.424 3.0685 0.516 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0465 0.576 1.3115 0.7035 ;
              RECT  1.0465 0.5585 1.177 0.7035 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.4665 0.523 0.774 ;
              RECT  0.4205 0.4665 0.523 0.6505 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.101 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.101 0.042 ;
        END
    END VSS
END SDFFRHQX2

MACRO CLKMX2X4
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.368 0.742 1.4105 1.0465 ;
              RECT  1.11 0.332 1.4105 0.3745 ;
              RECT  1.368 0.2755 1.4105 0.3745 ;
              RECT  1.078 0.742 1.4105 0.7845 ;
              RECT  1.11 0.6925 1.23 0.7845 ;
              RECT  1.11 0.2965 1.1525 0.7845 ;
              RECT  1.078 0.742 1.1205 1.0465 ;
              RECT  1.057 0.2965 1.1525 0.339 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.873 0.576 1.039 0.6325 ;
              RECT  0.834 0.6715 0.9295 0.781 ;
              RECT  0.873 0.576 0.9295 0.781 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.445 0.3815 0.799 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4525 0.643 0.537 0.6855 ;
              RECT  0.1835 0.8695 0.4945 0.912 ;
              RECT  0.4525 0.643 0.4945 0.912 ;
              RECT  0.1835 0.6925 0.24 0.912 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END CLKMX2X4

MACRO EDFFTRX2
    CLASS CORE ;
    SIZE 5.515 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.992 0.728 5.1015 0.7845 ;
              RECT  4.992 0.6925 5.052 0.7845 ;
              RECT  4.9955 0.3815 5.052 0.7845 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.7195 0.5585 4.907 0.6505 ;
              RECT  4.6845 0.7495 4.7765 0.806 ;
              RECT  4.7195 0.3815 4.7765 0.806 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.4085 0.7105 4.5005 0.767 ;
              RECT  4.444 0.449 4.5005 0.767 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8805 0.53 1.937 0.8835 ;
        END
    END RN
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9225 0.544 1.0465 0.5865 ;
              RECT  0.4985 0.7705 0.965 0.813 ;
              RECT  0.9225 0.544 0.965 0.813 ;
              RECT  0.4985 0.516 0.5405 0.813 ;
              RECT  0.449 0.7105 0.5405 0.767 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.424 0.3955 0.516 ;
              RECT  0.1835 0.424 0.24 0.622 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 5.515 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 5.515 0.042 ;
        END
    END VSS
END EDFFTRX2

MACRO CLKAND2X6
    CLASS CORE ;
    SIZE 1.9795 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.8875 0.608 1.93 0.9685 ;
              RECT  1.269 0.371 1.8915 0.4135 ;
              RECT  1.849 0.194 1.8915 0.4135 ;
              RECT  1.308 0.608 1.93 0.6505 ;
              RECT  1.739 0.5585 1.796 0.6505 ;
              RECT  1.739 0.371 1.7815 0.6505 ;
              RECT  1.598 0.608 1.64 0.9685 ;
              RECT  1.559 0.194 1.6015 0.4135 ;
              RECT  1.308 0.608 1.3505 0.9685 ;
              RECT  1.269 0.194 1.3115 0.4135 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3815 0.576 0.841 0.6325 ;
              RECT  0.7565 0.555 0.841 0.6325 ;
              RECT  0.3815 0.555 0.4665 0.6325 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.0425 0.4415 1.085 0.5265 ;
              RECT  0.166 0.4415 1.085 0.484 ;
              RECT  0.1235 0.456 0.258 0.4985 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.9795 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.9795 0.042 ;
        END
    END VSS
END CLKAND2X6

MACRO OA21X2
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.905 0.403 1.057 0.445 ;
              RECT  0.8905 0.424 0.9475 0.516 ;
              RECT  0.8485 0.4735 0.8905 1.0285 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.3955 0.24 0.7495 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.555 0.4985 0.6115 ;
              RECT  0.4415 0.417 0.4985 0.6115 ;
              RECT  0.325 0.555 0.3815 0.654 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.1555 0.6645 0.509 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END OA21X2

MACRO OAI31X2
    CLASS CORE ;
    SIZE 1.5555 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.202 0.385 1.3255 0.4275 ;
              RECT  1.202 0.385 1.2445 0.7845 ;
              RECT  1.17 0.742 1.2125 1.0145 ;
              RECT  0.643 0.8375 1.2125 0.88 ;
              RECT  1.032 0.742 1.2125 0.88 ;
              RECT  1.032 0.6925 1.0885 0.88 ;
              RECT  0.643 0.8375 0.6855 0.9225 ;
        END
    END Y
    PIN A2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.668 0.647 0.919 0.7035 ;
              RECT  0.629 0.7105 0.8235 0.767 ;
              RECT  0.668 0.647 0.8235 0.767 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.35 0.5335 0.873 0.576 ;
              RECT  0.4665 0.5335 0.523 0.6505 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.9895 0.424 1.0885 0.5795 ;
              RECT  0.2365 0.4205 1.032 0.463 ;
              RECT  0.2365 0.4205 0.279 0.562 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.315 0.4985 1.3715 0.852 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.5555 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.5555 0.042 ;
        END
    END VSS
END OAI31X2

MACRO EDFFHQX1
    CLASS CORE ;
    SIZE 3.5355 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.1635 0.5585 2.2485 0.7705 ;
              RECT  2.192 0.378 2.2485 0.7705 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.2205 0.4415 3.369 0.5055 ;
              RECT  2.959 0.4415 3.369 0.484 ;
              RECT  3.0405 0.2155 3.0825 0.484 ;
              RECT  2.7115 0.2155 3.0825 0.258 ;
              RECT  2.959 0.4415 3.0015 0.5265 ;
              RECT  2.7115 0.2155 2.754 0.6395 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.0935 0.576 3.3725 0.661 ;
              RECT  3.0935 0.555 3.15 0.6855 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.516 0.24 0.8695 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.5355 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.5355 0.042 ;
        END
    END VSS
END EDFFHQX1

MACRO SDFFSRX2
    CLASS CORE ;
    SIZE 6.6465 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  6.109 0.403 6.194 0.445 ;
              RECT  6.109 0.403 6.1515 0.9225 ;
              RECT  5.982 0.4735 6.1515 0.516 ;
              RECT  5.982 0.424 6.0385 0.516 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.7415 0.3815 5.798 0.9225 ;
              RECT  5.699 0.6925 5.798 0.7845 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  5.3985 0.6715 5.5575 0.767 ;
              RECT  5.3985 0.516 5.455 0.767 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.266 0.477 2.5525 0.5335 ;
              RECT  2.266 0.4415 2.379 0.5655 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.371 1.23 0.7245 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.032 0.424 1.0885 0.516 ;
              RECT  0.905 0.424 1.0885 0.4805 ;
              RECT  0.905 0.424 0.9615 0.615 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4275 0.5055 0.484 0.7565 ;
              RECT  0.325 0.5055 0.484 0.6505 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7915 0.1625 0.834 0.728 ;
              RECT  0.463 0.1625 0.834 0.205 ;
              RECT  0.523 0.3955 0.608 0.438 ;
              RECT  0.1975 0.392 0.548 0.4345 ;
              RECT  0.463 0.1625 0.5055 0.4345 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 6.6465 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 6.6465 0.042 ;
        END
    END VSS
END SDFFSRX2

MACRO OA22X4
    CLASS CORE ;
    SIZE 1.697 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8765 0.742 1.513 0.7845 ;
              RECT  1.375 0.6925 1.513 0.7845 ;
              RECT  1.375 0.2895 1.4175 0.7845 ;
              RECT  1.103 0.325 1.4175 0.3675 ;
              RECT  1.1665 0.742 1.209 1.018 ;
              RECT  1.0535 0.311 1.138 0.3535 ;
              RECT  0.8765 0.742 0.919 1.018 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.6925 0.806 0.8625 ;
              RECT  0.707 0.5515 0.7635 0.7495 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.622 0.3955 0.8485 ;
              RECT  0.339 0.509 0.3955 0.8485 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.509 0.24 0.8625 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.509 0.523 0.8625 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.697 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.697 0.042 ;
        END
    END VSS
END OA22X4

MACRO CLKAND2X3
    CLASS CORE ;
    SIZE 1.2725 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1065 0.668 1.149 0.9435 ;
              RECT  0.795 0.35 1.1065 0.392 ;
              RECT  1.064 0.293 1.1065 0.392 ;
              RECT  0.8165 0.668 1.149 0.7105 ;
              RECT  1.032 0.35 1.0885 0.7105 ;
              RECT  0.8165 0.668 0.859 0.9435 ;
              RECT  0.753 0.3145 0.8375 0.357 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1625 0.569 0.403 0.654 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.152 0.4415 0.569 0.4985 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 1.2725 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 1.2725 0.042 ;
        END
    END VSS
END CLKAND2X3

MACRO EDFFX2
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.309 0.357 3.4045 0.3995 ;
              RECT  3.309 0.357 3.3515 0.958 ;
              RECT  3.295 0.424 3.3515 0.516 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.9945 0.4415 3.0865 0.4985 ;
              RECT  2.9945 0.357 3.072 0.4985 ;
              RECT  2.9945 0.357 3.037 0.958 ;
              RECT  2.9875 0.357 3.072 0.3995 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.7115 0.576 2.8035 0.6325 ;
              RECT  2.7115 0.548 2.7965 0.6325 ;
              RECT  1.983 0.8835 2.7715 0.926 ;
              RECT  2.729 0.548 2.7715 0.926 ;
              RECT  2.1315 0.47 2.174 0.926 ;
              RECT  2.0895 0.47 2.174 0.5125 ;
              RECT  1.941 1.0075 2.0255 1.05 ;
              RECT  1.983 0.8835 2.0255 1.05 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4005 0.4525 2.5275 0.509 ;
              RECT  2.4465 0.4525 2.503 0.735 ;
              RECT  2.4005 0.4525 2.503 0.5125 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1625 0.548 0.286 0.6325 ;
              RECT  0.2295 0.438 0.286 0.6325 ;
              RECT  0.166 0.548 0.2225 0.7245 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END EDFFX2

MACRO DLY3X1
    CLASS CORE ;
    SIZE 3.394 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.001 0.576 2.0435 0.912 ;
              RECT  1.863 0.576 2.0435 0.6325 ;
              RECT  1.863 0.3815 1.9055 0.6325 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.1735 0.5585 1.368 0.753 ;
              RECT  1.2405 0.537 1.368 0.753 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.394 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.394 0.042 ;
        END
    END VSS
END DLY3X1

MACRO OAI222X4
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5775 0.5585 3.6345 0.6505 ;
              RECT  3.581 0.378 3.6235 0.6505 ;
              RECT  0.548 0.8165 3.62 0.859 ;
              RECT  3.5775 0.4345 3.62 0.859 ;
              RECT  2.7115 0.4345 3.6235 0.477 ;
              RECT  3.2915 0.378 3.334 0.477 ;
              RECT  3.2735 0.8165 3.316 0.9015 ;
              RECT  3.0015 0.378 3.044 0.477 ;
              RECT  2.8315 0.8165 2.874 0.9015 ;
              RECT  2.7115 0.378 2.754 0.477 ;
              RECT  2.2765 0.8165 2.319 0.9015 ;
              RECT  1.672 0.8165 1.7145 0.9015 ;
              RECT  1.0215 0.8165 1.064 0.9015 ;
              RECT  0.548 0.8165 0.59 0.9015 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.2155 0.7035 1.23 0.7455 ;
              RECT  1.1735 0.5585 1.23 0.7455 ;
              RECT  0.753 0.661 0.8375 0.7455 ;
              RECT  0.2155 0.661 0.258 0.7455 ;
        END
    END A0
    PIN C0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.729 0.7035 3.4825 0.7455 ;
              RECT  3.44 0.6325 3.4825 0.7455 ;
              RECT  3.0755 0.661 3.1605 0.7455 ;
              RECT  2.729 0.5585 2.786 0.7455 ;
              RECT  2.6375 0.59 2.786 0.6325 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.4465 0.5585 2.503 0.6505 ;
              RECT  1.474 0.7035 2.489 0.7455 ;
              RECT  2.4465 0.5585 2.489 0.7455 ;
              RECT  1.8985 0.661 1.983 0.7455 ;
              RECT  1.474 0.6325 1.5165 0.7455 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4735 0.548 1.039 0.59 ;
              RECT  0.59 0.548 0.682 0.6325 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.277 0.548 3.369 0.6325 ;
              RECT  2.8565 0.548 3.369 0.59 ;
        END
    END C1
    PIN B1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  1.7215 0.548 2.2485 0.59 ;
              RECT  1.7215 0.548 1.8275 0.6325 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END OAI222X4

MACRO INVX2
    CLASS CORE ;
    SIZE 0.424 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.3285 0.3815 0.378 0.502 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.049 0.424 0.1235 0.5655 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.424 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.424 0.042 ;
        END
    END VSS
END INVX2

MACRO TLATNSRXL
    CLASS CORE ;
    SIZE 3.2525 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN QN
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.689 0.728 0.7455 0.8305 ;
              RECT  0.608 0.385 0.7455 0.4415 ;
              RECT  0.689 0.357 0.7455 0.4415 ;
              RECT  0.608 0.728 0.7455 0.7845 ;
              RECT  0.608 0.385 0.6645 0.7845 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.173 0.3815 0.2295 0.721 ;
              RECT  0.042 0.424 0.2295 0.516 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.012 0.5865 3.118 0.7845 ;
              RECT  3.012 0.5865 3.0685 0.8905 ;
        END
    END GN
    PIN RN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.588 0.608 2.9415 0.6505 ;
              RECT  2.588 0.5585 2.6795 0.6505 ;
              RECT  2.6375 0.2435 2.6795 0.6505 ;
              RECT  1.301 0.2435 2.6795 0.286 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.082 0.47 2.2485 0.6505 ;
              RECT  2.082 0.47 2.1385 0.714 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.8305 0.8445 0.965 0.9015 ;
              RECT  0.9085 0.6255 0.965 0.9015 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.2525 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.2525 0.042 ;
        END
    END VSS
END TLATNSRXL

MACRO MXI2XL
    CLASS CORE ;
    SIZE 0.9895 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.385 0.852 0.4275 0.9365 ;
              RECT  0.1975 0.852 0.4275 0.894 ;
              RECT  0.1975 0.339 0.3675 0.3815 ;
              RECT  0.1975 0.339 0.24 0.894 ;
              RECT  0.1835 0.424 0.24 0.516 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7495 0.5655 0.806 0.7845 ;
              RECT  0.463 0.5655 0.806 0.622 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.544 0.6925 0.6785 0.8485 ;
        END
    END B
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.0705 0.5935 0.127 0.8485 ;
              RECT  0.042 0.523 0.0985 0.6505 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.9895 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.9895 0.042 ;
        END
    END VSS
END MXI2XL

MACRO NAND4XL
    CLASS CORE ;
    SIZE 0.8485 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Y
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.258 0.675 0.806 0.7175 ;
              RECT  0.7635 0.2895 0.806 0.7175 ;
              RECT  0.7495 0.2895 0.806 0.449 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.251 0.24 0.6045 ;
        END
    END A
    PIN B
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.325 0.251 0.3815 0.6045 ;
        END
    END B
    PIN C
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.4665 0.251 0.523 0.6045 ;
        END
    END C
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.608 0.251 0.6645 0.6045 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 0.8485 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 0.8485 0.042 ;
        END
    END VSS
END NAND4XL

MACRO DFFHQX8
    CLASS CORE ;
    SIZE 3.818 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.5635 0.4735 3.6695 0.6645 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.4365 0.555 3.493 0.6645 ;
              RECT  3.2735 0.555 3.493 0.6505 ;
              RECT  3.2735 0.4735 3.33 0.6505 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.926 0.3815 0.9685 0.951 ;
              RECT  0.346 0.424 0.9685 0.4665 ;
              RECT  0.636 0.3815 0.6785 0.951 ;
              RECT  0.346 0.3815 0.3885 0.951 ;
              RECT  0.042 0.4735 0.3885 0.516 ;
              RECT  0.0565 0.3815 0.0985 0.951 ;
              RECT  0.042 0.424 0.0985 0.516 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 3.818 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 3.818 0.042 ;
        END
    END VSS
END DFFHQX8

MACRO EDFFHQX4
    CLASS CORE ;
    SIZE 4.384 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN Q
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.6725 0.403 2.7575 0.445 ;
              RECT  2.1775 0.53 2.715 0.5725 ;
              RECT  2.6725 0.403 2.715 0.5725 ;
              RECT  2.2415 0.795 2.6335 0.8375 ;
              RECT  2.2375 0.7105 2.28 0.82 ;
              RECT  2.146 0.7105 2.28 0.767 ;
              RECT  2.1775 0.403 2.22 0.767 ;
              RECT  2.135 0.403 2.22 0.445 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  4.1255 0.4415 4.2175 0.4985 ;
              RECT  4.1255 0.3425 4.168 0.4985 ;
              RECT  3.7475 0.3425 4.168 0.385 ;
              RECT  3.705 0.4415 3.79 0.484 ;
              RECT  3.7475 0.173 3.79 0.484 ;
              RECT  3.4785 0.173 3.79 0.2155 ;
              RECT  3.4785 0.173 3.521 0.647 ;
        END
    END E
    PIN D
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  3.8605 0.5585 4.055 0.6715 ;
              RECT  3.9985 0.456 4.055 0.6715 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.1835 0.5725 0.24 0.926 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 4.384 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 4.384 0.042 ;
        END
    END VSS
END EDFFHQX4

MACRO TLATNCAX4
    CLASS CORE ;
    SIZE 2.5455 BY 1.209 ;
    SYMMETRY X Y ;
    SITE CoreSiteDie1 ;
    PIN ECK
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.7635 0.6575 0.8485 0.7 ;
              RECT  0.7455 0.3885 0.8305 0.431 ;
              RECT  0.4525 0.636 0.806 0.6785 ;
              RECT  0.4665 0.403 0.781 0.445 ;
              RECT  0.4665 0.5585 0.523 0.6785 ;
              RECT  0.4665 0.3605 0.509 0.6785 ;
              RECT  0.4525 0.636 0.4945 0.721 ;
        END
    END ECK
    PIN E
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  2.0855 0.5515 2.298 0.6325 ;
              RECT  2.0855 0.5515 2.1425 0.7495 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0.233 0.4595 0.3815 0.516 ;
              RECT  0.325 0.424 0.3815 0.516 ;
              RECT  0.233 0.4595 0.2895 0.6855 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 1.1665 2.5455 1.209 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT
            LAYER Metal1Die1 ;
              RECT  0 0 2.5455 0.042 ;
        END
    END VSS
END TLATNCAX4
END LIBRARY
