VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.1 ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.042 ;
END M1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
END M2

SITE site1
  CLASS CORE ;
  SIZE 50 BY 20 ;
END site1

MACRO BUF_X1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END BUF_X1

MACRO BUF_X2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END BUF_X2

MACRO INV_X1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ;
    DIRECTION OUTPUT ;
    PORT
        LAYER M1 ;
            RECT 40 15 45 20 ;
    END
 END ZN
 PIN A DIRECTION INPUT ;
    DIRECTION INPUT ;
    PORT
        LAYER M1 ;
            RECT 5 5 10 10 ;
    END
 END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END INV_X1

MACRO AND2_X1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ;
     PORT
         LAYER M1 ;
             RECT 40 15 45 20 ;
     END
 END ZN
 PIN A1
    DIRECTION INPUT ;
    PORT
        LAYER M1 ;
            RECT 10 10 15 15 ;
    END
 END A1
 PIN A2 DIRECTION INPUT ; END A2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END AND2_X1

MACRO NOR2_X1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A1 DIRECTION INPUT ; END A1
 PIN A2 DIRECTION INPUT ; END A2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END NOR2_X1

MACRO DFF_X1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ;
      PORT
          LAYER M1 ;
              RECT 40 10 45 15 ;
      END
 END Q
 PIN D DIRECTION INPUT ;
     DIRECTION INPUT ;
     PORT
         LAYER M1 ;
             RECT 10 10 15 15 ;
     END
 END D
 PIN CK DIRECTION INPUT ;
     DIRECTION INPUT ;
     PORT
         LAYER M1 ;
             RECT 23 0 25 5 ;
     END
 END CK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END DFF_X1

END LIBRARY
