VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.1 ;

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.042 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.08 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
END metal2

LAYER metal3
  TYPE ROUTING ;
  SPACINGTABLE
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.88 ;
  CAPACITANCE CPERSQDIST 2.7745e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  SPACINGTABLE
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.14 ;
  CAPACITANCE CPERSQDIST 2.0743e-05 ;
  EDGECAPACITANCE 3.0908e-05 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  SPACINGTABLE
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.71 ;
  CAPACITANCE CPERSQDIST 1.3527e-05 ;
  EDGECAPACITANCE 2.3863e-06 ;
END metal5


SITE site1
  CLASS CORE ;
  SIZE 50 BY 20 ;
END site1

MACRO BUF_X1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END BUF_X1

MACRO BUF_X2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END BUF_X2

MACRO INV_X1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ;
    DIRECTION OUTPUT ;
    PORT
        LAYER metal1 ;
            RECT 40 15 45 20 ;
    END
 END ZN
 PIN A DIRECTION INPUT ;
    DIRECTION INPUT ;
    PORT
        LAYER metal1 ;
            RECT 5 5 10 10 ;
    END
 END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END INV_X1

MACRO AND2_X1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ;
     PORT
         LAYER metal1 ;
             RECT 40 15 45 20 ;
     END
 END ZN
 PIN A1
    DIRECTION INPUT ;
    PORT
        LAYER metal1 ;
            RECT 10 10 15 15 ;
    END
 END A1
 PIN A2 DIRECTION INPUT ; END A2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END AND2_X1

MACRO NOR2_X1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A1 DIRECTION INPUT ; END A1
 PIN A2 DIRECTION INPUT ; END A2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END NOR2_X1

MACRO DFF_X1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ;
      PORT
          LAYER metal1 ;
              RECT 40 10 45 15 ;
      END
 END Q
 PIN D DIRECTION INPUT ;
     DIRECTION INPUT ;
     PORT
         LAYER metal1 ;
             RECT 10 10 15 15 ;
     END
 END D
 PIN CK DIRECTION INPUT ;
     DIRECTION INPUT ;
     PORT
         LAYER metal1 ;
             RECT 23 0 25 5 ;
     END
 END CK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END DFF_X1

END LIBRARY
